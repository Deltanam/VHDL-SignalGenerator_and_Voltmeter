
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Triangle_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    STD_LOGIC_VECTOR(8 DOWNTO 0);                           
      duty_cycle     :  OUT   STD_LOGIC_VECTOR(8 DOWNTO 0)
		);
END Triangle_Lookup;

ARCHITECTURE behavior OF Triangle_Lookup IS

type array_1d is array (0 to 511) of integer;

constant triangle : array_1d := (				
(	0	)	,
(	2	)	,
(	4	)	,
(	6	)	,
(	8	)	,
(	10	)	,
(	12	)	,
(	14	)	,
(	16	)	,
(	18	)	,
(	20	)	,
(	22	)	,
(	24	)	,
(	26	)	,
(	28	)	,
(	30	)	,
(	32	)	,
(	34	)	,
(	36	)	,
(	38	)	,
(	40	)	,
(	42	)	,
(	44	)	,
(	46	)	,
(	48	)	,
(	50	)	,
(	52	)	,
(	54	)	,
(	56	)	,
(	58	)	,
(	60	)	,
(	62	)	,
(	64	)	,
(	66	)	,
(	68	)	,
(	70	)	,
(	72	)	,
(	74	)	,
(	76	)	,
(	78	)	,
(	80	)	,
(	82	)	,
(	84	)	,
(	86	)	,
(	88	)	,
(	90	)	,
(	92	)	,
(	94	)	,
(	96	)	,
(	98	)	,
(	100	)	,
(	102	)	,
(	104	)	,
(	106	)	,
(	108	)	,
(	110	)	,
(	112	)	,
(	114	)	,
(	116	)	,
(	118	)	,
(	120	)	,
(	122	)	,
(	124	)	,
(	126	)	,
(	128	)	,
(	130	)	,
(	132	)	,
(	134	)	,
(	136	)	,
(	138	)	,
(	140	)	,
(	142	)	,
(	144	)	,
(	146	)	,
(	148	)	,
(	150	)	,
(	152	)	,
(	154	)	,
(	156	)	,
(	158	)	,
(	160	)	,
(	162	)	,
(	164	)	,
(	166	)	,
(	168	)	,
(	170	)	,
(	172	)	,
(	174	)	,
(	176	)	,
(	178	)	,
(	180	)	,
(	182	)	,
(	184	)	,
(	186	)	,
(	188	)	,
(	190	)	,
(	192	)	,
(	194	)	,
(	196	)	,
(	198	)	,
(	200	)	,
(	202	)	,
(	204	)	,
(	206	)	,
(	208	)	,
(	210	)	,
(	212	)	,
(	214	)	,
(	216	)	,
(	218	)	,
(	220	)	,
(	222	)	,
(	224	)	,
(	226	)	,
(	228	)	,
(	230	)	,
(	232	)	,
(	234	)	,
(	236	)	,
(	238	)	,
(	240	)	,
(	242	)	,
(	244	)	,
(	246	)	,
(	248	)	,
(	250	)	,
(	252	)	,
(	254	)	,
(	256	)	,
(	258	)	,
(	260	)	,
(	262	)	,
(	264	)	,
(	266	)	,
(	268	)	,
(	270	)	,
(	272	)	,
(	274	)	,
(	276	)	,
(	278	)	,
(	280	)	,
(	282	)	,
(	284	)	,
(	286	)	,
(	288	)	,
(	290	)	,
(	292	)	,
(	294	)	,
(	296	)	,
(	298	)	,
(	300	)	,
(	302	)	,
(	304	)	,
(	306	)	,
(	308	)	,
(	310	)	,
(	312	)	,
(	314	)	,
(	316	)	,
(	318	)	,
(	320	)	,
(	322	)	,
(	324	)	,
(	326	)	,
(	328	)	,
(	330	)	,
(	332	)	,
(	334	)	,
(	336	)	,
(	338	)	,
(	340	)	,
(	342	)	,
(	344	)	,
(	346	)	,
(	348	)	,
(	350	)	,
(	352	)	,
(	354	)	,
(	356	)	,
(	358	)	,
(	360	)	,
(	362	)	,
(	364	)	,
(	366	)	,
(	368	)	,
(	370	)	,
(	372	)	,
(	374	)	,
(	376	)	,
(	378	)	,
(	380	)	,
(	382	)	,
(	384	)	,
(	386	)	,
(	388	)	,
(	390	)	,
(	392	)	,
(	394	)	,
(	396	)	,
(	398	)	,
(	400	)	,
(	402	)	,
(	404	)	,
(	406	)	,
(	408	)	,
(	410	)	,
(	412	)	,
(	414	)	,
(	416	)	,
(	418	)	,
(	420	)	,
(	422	)	,
(	424	)	,
(	426	)	,
(	428	)	,
(	430	)	,
(	432	)	,
(	434	)	,
(	436	)	,
(	438	)	,
(	440	)	,
(	442	)	,
(	444	)	,
(	446	)	,
(	448	)	,
(	450	)	,
(	452	)	,
(	454	)	,
(	456	)	,
(	458	)	,
(	460	)	,
(	462	)	,
(	464	)	,
(	466	)	,
(	468	)	,
(	470	)	,
(	472	)	,
(	474	)	,
(	476	)	,
(	478	)	,
(	480	)	,
(	482	)	,
(	484	)	,
(	486	)	,
(	488	)	,
(	490	)	,
(	492	)	,
(	494	)	,
(	496	)	,
(	498	)	,
(	500	)	,
(	502	)	,
(	504	)	,
(	506	)	,
(	508	)	,
(	510	)	,
(	511	)	,
(	509	)	,
(	507	)	,
(	505	)	,
(	503	)	,
(	501	)	,
(	499	)	,
(	497	)	,
(	495	)	,
(	493	)	,
(	491	)	,
(	489	)	,
(	487	)	,
(	485	)	,
(	483	)	,
(	481	)	,
(	479	)	,
(	477	)	,
(	475	)	,
(	473	)	,
(	471	)	,
(	469	)	,
(	467	)	,
(	465	)	,
(	463	)	,
(	461	)	,
(	459	)	,
(	457	)	,
(	455	)	,
(	453	)	,
(	451	)	,
(	449	)	,
(	447	)	,
(	445	)	,
(	443	)	,
(	441	)	,
(	439	)	,
(	437	)	,
(	435	)	,
(	433	)	,
(	431	)	,
(	429	)	,
(	427	)	,
(	425	)	,
(	423	)	,
(	421	)	,
(	419	)	,
(	417	)	,
(	415	)	,
(	413	)	,
(	411	)	,
(	409	)	,
(	407	)	,
(	405	)	,
(	403	)	,
(	401	)	,
(	399	)	,
(	397	)	,
(	395	)	,
(	393	)	,
(	391	)	,
(	389	)	,
(	387	)	,
(	385	)	,
(	383	)	,
(	381	)	,
(	379	)	,
(	377	)	,
(	375	)	,
(	373	)	,
(	371	)	,
(	369	)	,
(	367	)	,
(	365	)	,
(	363	)	,
(	361	)	,
(	359	)	,
(	357	)	,
(	355	)	,
(	353	)	,
(	351	)	,
(	349	)	,
(	347	)	,
(	345	)	,
(	343	)	,
(	341	)	,
(	339	)	,
(	337	)	,
(	335	)	,
(	333	)	,
(	331	)	,
(	329	)	,
(	327	)	,
(	325	)	,
(	323	)	,
(	321	)	,
(	319	)	,
(	317	)	,
(	315	)	,
(	313	)	,
(	311	)	,
(	309	)	,
(	307	)	,
(	305	)	,
(	303	)	,
(	301	)	,
(	299	)	,
(	297	)	,
(	295	)	,
(	293	)	,
(	291	)	,
(	289	)	,
(	287	)	,
(	285	)	,
(	283	)	,
(	281	)	,
(	279	)	,
(	277	)	,
(	275	)	,
(	273	)	,
(	271	)	,
(	269	)	,
(	267	)	,
(	265	)	,
(	263	)	,
(	261	)	,
(	259	)	,
(	257	)	,
(	255	)	,
(	253	)	,
(	251	)	,
(	249	)	,
(	247	)	,
(	245	)	,
(	243	)	,
(	241	)	,
(	239	)	,
(	237	)	,
(	235	)	,
(	233	)	,
(	231	)	,
(	229	)	,
(	227	)	,
(	225	)	,
(	223	)	,
(	221	)	,
(	219	)	,
(	217	)	,
(	215	)	,
(	213	)	,
(	211	)	,
(	209	)	,
(	207	)	,
(	205	)	,
(	203	)	,
(	201	)	,
(	199	)	,
(	197	)	,
(	195	)	,
(	193	)	,
(	191	)	,
(	189	)	,
(	187	)	,
(	185	)	,
(	183	)	,
(	181	)	,
(	179	)	,
(	177	)	,
(	175	)	,
(	173	)	,
(	171	)	,
(	169	)	,
(	167	)	,
(	165	)	,
(	163	)	,
(	161	)	,
(	159	)	,
(	157	)	,
(	155	)	,
(	153	)	,
(	151	)	,
(	149	)	,
(	147	)	,
(	145	)	,
(	143	)	,
(	141	)	,
(	139	)	,
(	137	)	,
(	135	)	,
(	133	)	,
(	131	)	,
(	129	)	,
(	127	)	,
(	125	)	,
(	123	)	,
(	121	)	,
(	119	)	,
(	117	)	,
(	115	)	,
(	113	)	,
(	111	)	,
(	109	)	,
(	107	)	,
(	105	)	,
(	103	)	,
(	101	)	,
(	99	)	,
(	97	)	,
(	95	)	,
(	93	)	,
(	91	)	,
(	89	)	,
(	87	)	,
(	85	)	,
(	83	)	,
(	81	)	,
(	79	)	,
(	77	)	,
(	75	)	,
(	73	)	,
(	71	)	,
(	69	)	,
(	67	)	,
(	65	)	,
(	63	)	,
(	61	)	,
(	59	)	,
(	57	)	,
(	55	)	,
(	53	)	,
(	51	)	,
(	49	)	,
(	47	)	,
(	45	)	,
(	43	)	,
(	41	)	,
(	39	)	,
(	37	)	,
(	35	)	,
(	33	)	,
(	31	)	,
(	29	)	,
(	27	)	,
(	25	)	,
(	23	)	,
(	21	)	,
(	19	)	,
(	17	)	,
(	15	)	,
(	13	)	,
(	11	)	,
(	9	)	,
(	7	)	,
(	5	)	,
(	3	)	,
(	1	)


);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	
	duty_cycle <= std_logic_vector(to_unsigned(triangle(to_integer(unsigned(index))),duty_cycle'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
