
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY BuzzFreq_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    integer;                           
      Divisor     :  OUT   natural
		);
END BuzzFreq_Lookup;

ARCHITECTURE behavior OF BuzzFreq_Lookup IS

type array_1d is array (0 to 4095) of natural;

constant Divisors : array_1d := (				

(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	1286008	)	,
(	1262626	)	,
(	1240079	)	,
(	1218324	)	,
(	1197318	)	,
(	1177024	)	,
(	1157407	)	,
(	1138434	)	,
(	1120072	)	,
(	1102293	)	,
(	1085069	)	,
(	1068376	)	,
(	1052189	)	,
(	1036484	)	,
(	1021242	)	,
(	1006441	)	,
(	992063	)	,
(	978091	)	,
(	964506	)	,
(	951294	)	,
(	938438	)	,
(	925926	)	,
(	913743	)	,
(	901876	)	,
(	890313	)	,
(	879044	)	,
(	868056	)	,
(	857339	)	,
(	846883	)	,
(	836680	)	,
(	826720	)	,
(	816993	)	,
(	807494	)	,
(	798212	)	,
(	789141	)	,
(	780275	)	,
(	771605	)	,
(	763126	)	,
(	754831	)	,
(	746714	)	,
(	738771	)	,
(	730994	)	,
(	723380	)	,
(	715922	)	,
(	708617	)	,
(	701459	)	,
(	694444	)	,
(	687569	)	,
(	680828	)	,
(	674218	)	,
(	667735	)	,
(	661376	)	,
(	655136	)	,
(	649013	)	,
(	643004	)	,
(	637105	)	,
(	631313	)	,
(	625626	)	,
(	620040	)	,
(	614553	)	,
(	609162	)	,
(	603865	)	,
(	598659	)	,
(	593542	)	,
(	588512	)	,
(	583567	)	,
(	578704	)	,
(	573921	)	,
(	569217	)	,
(	564589	)	,
(	560036	)	,
(	555556	)	,
(	551146	)	,
(	546807	)	,
(	542535	)	,
(	538329	)	,
(	534188	)	,
(	530110	)	,
(	526094	)	,
(	522139	)	,
(	518242	)	,
(	514403	)	,
(	510621	)	,
(	506894	)	,
(	503221	)	,
(	499600	)	,
(	496032	)	,
(	492514	)	,
(	489045	)	,
(	485625	)	,
(	482253	)	,
(	478927	)	,
(	475647	)	,
(	472411	)	,
(	469219	)	,
(	466070	)	,
(	462963	)	,
(	459897	)	,
(	456871	)	,
(	453885	)	,
(	450938	)	,
(	448029	)	,
(	445157	)	,
(	442321	)	,
(	439522	)	,
(	436758	)	,
(	434028	)	,
(	431332	)	,
(	428669	)	,
(	426040	)	,
(	423442	)	,
(	420875	)	,
(	418340	)	,
(	415835	)	,
(	413360	)	,
(	410914	)	,
(	408497	)	,
(	406108	)	,
(	403747	)	,
(	401413	)	,
(	399106	)	,
(	396825	)	,
(	394571	)	,
(	392341	)	,
(	390137	)	,
(	387958	)	,
(	385802	)	,
(	383671	)	,
(	381563	)	,
(	379478	)	,
(	377415	)	,
(	375375	)	,
(	373357	)	,
(	371361	)	,
(	369385	)	,
(	367431	)	,
(	365497	)	,
(	363583	)	,
(	361690	)	,
(	359816	)	,
(	357961	)	,
(	356125	)	,
(	354308	)	,
(	352510	)	,
(	350730	)	,
(	348967	)	,
(	347222	)	,
(	345495	)	,
(	343784	)	,
(	342091	)	,
(	340414	)	,
(	338753	)	,
(	337109	)	,
(	335480	)	,
(	333868	)	,
(	332270	)	,
(	330688	)	,
(	329121	)	,
(	327568	)	,
(	326030	)	,
(	324507	)	,
(	322997	)	,
(	321502	)	,
(	320020	)	,
(	318552	)	,
(	317098	)	,
(	315657	)	,
(	314228	)	,
(	312813	)	,
(	311410	)	,
(	310020	)	,
(	308642	)	,
(	307276	)	,
(	305923	)	,
(	304581	)	,
(	303251	)	,
(	301932	)	,
(	300625	)	,
(	299330	)	,
(	298045	)	,
(	296771	)	,
(	295508	)	,
(	294256	)	,
(	293015	)	,
(	291783	)	,
(	290563	)	,
(	289352	)	,
(	288151	)	,
(	286961	)	,
(	285780	)	,
(	284608	)	,
(	283447	)	,
(	282294	)	,
(	281152	)	,
(	280018	)	,
(	278893	)	,
(	277778	)	,
(	276671	)	,
(	275573	)	,
(	274484	)	,
(	273403	)	,
(	272331	)	,
(	271267	)	,
(	270212	)	,
(	269165	)	,
(	268125	)	,
(	267094	)	,
(	266071	)	,
(	265055	)	,
(	264047	)	,
(	263047	)	,
(	262055	)	,
(	261069	)	,
(	260092	)	,
(	259121	)	,
(	258158	)	,
(	257202	)	,
(	256253	)	,
(	255310	)	,
(	254375	)	,
(	253447	)	,
(	252525	)	,
(	251610	)	,
(	250702	)	,
(	249800	)	,
(	248905	)	,
(	248016	)	,
(	247133	)	,
(	246257	)	,
(	245387	)	,
(	244523	)	,
(	243665	)	,
(	242813	)	,
(	241967	)	,
(	241127	)	,
(	240292	)	,
(	239464	)	,
(	238641	)	,
(	237823	)	,
(	237012	)	,
(	236206	)	,
(	235405	)	,
(	234610	)	,
(	233820	)	,
(	233035	)	,
(	232256	)	,
(	231481	)	,
(	230712	)	,
(	229948	)	,
(	229190	)	,
(	228436	)	,
(	227687	)	,
(	226943	)	,
(	226203	)	,
(	225469	)	,
(	224739	)	,
(	224014	)	,
(	223294	)	,
(	222578	)	,
(	221867	)	,
(	221161	)	,
(	220459	)	,
(	219761	)	,
(	219068	)	,
(	218379	)	,
(	217694	)	,
(	217014	)	,
(	216338	)	,
(	215666	)	,
(	214998	)	,
(	214335	)	,
(	213675	)	,
(	213020	)	,
(	212368	)	,
(	211721	)	,
(	211077	)	,
(	210438	)	,
(	209802	)	,
(	209170	)	,
(	208542	)	,
(	207917	)	,
(	207297	)	,
(	206680	)	,
(	206067	)	,
(	205457	)	,
(	204851	)	,
(	204248	)	,
(	203649	)	,
(	203054	)	,
(	202462	)	,
(	201873	)	,
(	201288	)	,
(	200706	)	,
(	200128	)	,
(	199553	)	,
(	198981	)	,
(	198413	)	,
(	197847	)	,
(	197285	)	,
(	196726	)	,
(	196171	)	,
(	195618	)	,
(	195069	)	,
(	194522	)	,
(	193979	)	,
(	193439	)	,
(	192901	)	,
(	192367	)	,
(	191835	)	,
(	191307	)	,
(	190781	)	,
(	190259	)	,
(	189739	)	,
(	189222	)	,
(	188708	)	,
(	188196	)	,
(	187688	)	,
(	187182	)	,
(	186679	)	,
(	186178	)	,
(	185680	)	,
(	185185	)	,
(	184693	)	,
(	184203	)	,
(	183715	)	,
(	183231	)	,
(	182749	)	,
(	182269	)	,
(	181792	)	,
(	181317	)	,
(	180845	)	,
(	180375	)	,
(	179908	)	,
(	179443	)	,
(	178981	)	,
(	178520	)	,
(	178063	)	,
(	177607	)	,
(	177154	)	,
(	176703	)	,
(	176255	)	,
(	175809	)	,
(	175365	)	,
(	174923	)	,
(	174484	)	,
(	174046	)	,
(	173611	)	,
(	173178	)	,
(	172747	)	,
(	172319	)	,
(	171892	)	,
(	171468	)	,
(	171045	)	,
(	170625	)	,
(	170207	)	,
(	169791	)	,
(	169377	)	,
(	168965	)	,
(	168554	)	,
(	168146	)	,
(	167740	)	,
(	167336	)	,
(	166934	)	,
(	166533	)	,
(	166135	)	,
(	165739	)	,
(	165344	)	,
(	164951	)	,
(	164560	)	,
(	164171	)	,
(	163784	)	,
(	163399	)	,
(	163015	)	,
(	162633	)	,
(	162253	)	,
(	161875	)	,
(	161499	)	,
(	161124	)	,
(	160751	)	,
(	160380	)	,
(	160010	)	,
(	159642	)	,
(	159276	)	,
(	158912	)	,
(	158549	)	,
(	158188	)	,
(	157828	)	,
(	157470	)	,
(	157114	)	,
(	156759	)	,
(	156406	)	,
(	156055	)	,
(	155705	)	,
(	155357	)	,
(	155010	)	,
(	154665	)	,
(	154321	)	,
(	153979	)	,
(	153638	)	,
(	153299	)	,
(	152961	)	,
(	152625	)	,
(	152290	)	,
(	151957	)	,
(	151625	)	,
(	151295	)	,
(	150966	)	,
(	150639	)	,
(	150313	)	,
(	149988	)	,
(	149665	)	,
(	149343	)	,
(	149022	)	,
(	148703	)	,
(	148386	)	,
(	148069	)	,
(	147754	)	,
(	147440	)	,
(	147128	)	,
(	146817	)	,
(	146507	)	,
(	146199	)	,
(	145892	)	,
(	145586	)	,
(	145281	)	,
(	144978	)	,
(	144676	)	,
(	144375	)	,
(	144076	)	,
(	143777	)	,
(	143480	)	,
(	143184	)	,
(	142890	)	,
(	142596	)	,
(	142304	)	,
(	142013	)	,
(	141723	)	,
(	141435	)	,
(	141147	)	,
(	140861	)	,
(	140576	)	,
(	140292	)	,
(	140009	)	,
(	139727	)	,
(	139447	)	,
(	139167	)	,
(	138889	)	,
(	138612	)	,
(	138336	)	,
(	138061	)	,
(	137787	)	,
(	137514	)	,
(	137242	)	,
(	136971	)	,
(	136702	)	,
(	136433	)	,
(	136166	)	,
(	135899	)	,
(	135634	)	,
(	135369	)	,
(	135106	)	,
(	134844	)	,
(	134582	)	,
(	134322	)	,
(	134063	)	,
(	133804	)	,
(	133547	)	,
(	133291	)	,
(	133035	)	,
(	132781	)	,
(	132528	)	,
(	132275	)	,
(	132024	)	,
(	131773	)	,
(	131524	)	,
(	131275	)	,
(	131027	)	,
(	130780	)	,
(	130535	)	,
(	130290	)	,
(	130046	)	,
(	129803	)	,
(	129561	)	,
(	129319	)	,
(	129079	)	,
(	128839	)	,
(	128601	)	,
(	128363	)	,
(	128126	)	,
(	127890	)	,
(	127655	)	,
(	127421	)	,
(	127188	)	,
(	126955	)	,
(	126723	)	,
(	126493	)	,
(	126263	)	,
(	126033	)	,
(	125805	)	,
(	125578	)	,
(	125351	)	,
(	125125	)	,
(	124900	)	,
(	124676	)	,
(	124452	)	,
(	124230	)	,
(	124008	)	,
(	123787	)	,
(	123567	)	,
(	123347	)	,
(	123128	)	,
(	122911	)	,
(	122693	)	,
(	122477	)	,
(	122261	)	,
(	122046	)	,
(	121832	)	,
(	121619	)	,
(	121406	)	,
(	121194	)	,
(	120983	)	,
(	120773	)	,
(	120563	)	,
(	120354	)	,
(	120146	)	,
(	119939	)	,
(	119732	)	,
(	119526	)	,
(	119320	)	,
(	119116	)	,
(	118912	)	,
(	118708	)	,
(	118506	)	,
(	118304	)	,
(	118103	)	,
(	117902	)	,
(	117702	)	,
(	117503	)	,
(	117305	)	,
(	117107	)	,
(	116910	)	,
(	116713	)	,
(	116518	)	,
(	116322	)	,
(	116128	)	,
(	115934	)	,
(	115741	)	,
(	115548	)	,
(	115356	)	,
(	115165	)	,
(	114974	)	,
(	114784	)	,
(	114595	)	,
(	114406	)	,
(	114218	)	,
(	114030	)	,
(	113843	)	,
(	113657	)	,
(	113471	)	,
(	113286	)	,
(	113102	)	,
(	112918	)	,
(	112734	)	,
(	112552	)	,
(	112370	)	,
(	112188	)	,
(	112007	)	,
(	111827	)	,
(	111647	)	,
(	111468	)	,
(	111289	)	,
(	111111	)	,
(	110934	)	,
(	110757	)	,
(	110580	)	,
(	110405	)	,
(	110229	)	,
(	110055	)	,
(	109880	)	,
(	109707	)	,
(	109534	)	,
(	109361	)	,
(	109189	)	,
(	109018	)	,
(	108847	)	,
(	108677	)	,
(	108507	)	,
(	108338	)	,
(	108169	)	,
(	108001	)	,
(	107833	)	,
(	107666	)	,
(	107499	)	,
(	107333	)	,
(	107167	)	,
(	107002	)	,
(	106838	)	,
(	106673	)	,
(	106510	)	,
(	106347	)	,
(	106184	)	,
(	106022	)	,
(	105860	)	,
(	105699	)	,
(	105539	)	,
(	105379	)	,
(	105219	)	,
(	105060	)	,
(	104901	)	,
(	104743	)	,
(	104585	)	,
(	104428	)	,
(	104271	)	,
(	104115	)	,
(	103959	)	,
(	103803	)	,
(	103648	)	,
(	103494	)	,
(	103340	)	,
(	103186	)	,
(	103033	)	,
(	102881	)	,
(	102728	)	,
(	102577	)	,
(	102425	)	,
(	102275	)	,
(	102124	)	,
(	101974	)	,
(	101825	)	,
(	101676	)	,
(	101527	)	,
(	101379	)	,
(	101231	)	,
(	101084	)	,
(	100937	)	,
(	100790	)	,
(	100644	)	,
(	100498	)	,
(	100353	)	,
(	100208	)	,
(	100064	)	,
(	99920	)	,
(	99777	)	,
(	99633	)	,
(	99491	)	,
(	99348	)	,
(	99206	)	,
(	99065	)	,
(	98924	)	,
(	98783	)	,
(	98643	)	,
(	98503	)	,
(	98363	)	,
(	98224	)	,
(	98085	)	,
(	97947	)	,
(	97809	)	,
(	97672	)	,
(	97534	)	,
(	97398	)	,
(	97261	)	,
(	97125	)	,
(	96989	)	,
(	96854	)	,
(	96719	)	,
(	96585	)	,
(	96451	)	,
(	96317	)	,
(	96183	)	,
(	96050	)	,
(	95918	)	,
(	95785	)	,
(	95654	)	,
(	95522	)	,
(	95391	)	,
(	95260	)	,
(	95129	)	,
(	94999	)	,
(	94869	)	,
(	94740	)	,
(	94611	)	,
(	94482	)	,
(	94354	)	,
(	94226	)	,
(	94098	)	,
(	93971	)	,
(	93844	)	,
(	93717	)	,
(	93591	)	,
(	93465	)	,
(	93339	)	,
(	93214	)	,
(	93089	)	,
(	92964	)	,
(	92840	)	,
(	92716	)	,
(	92593	)	,
(	92469	)	,
(	92346	)	,
(	92224	)	,
(	92101	)	,
(	91979	)	,
(	91858	)	,
(	91736	)	,
(	91615	)	,
(	91495	)	,
(	91374	)	,
(	91254	)	,
(	91134	)	,
(	91015	)	,
(	90896	)	,
(	90777	)	,
(	90659	)	,
(	90540	)	,
(	90422	)	,
(	90305	)	,
(	90188	)	,
(	90071	)	,
(	89954	)	,
(	89838	)	,
(	89722	)	,
(	89606	)	,
(	89490	)	,
(	89375	)	,
(	89260	)	,
(	89146	)	,
(	89031	)	,
(	88917	)	,
(	88804	)	,
(	88690	)	,
(	88577	)	,
(	88464	)	,
(	88352	)	,
(	88239	)	,
(	88127	)	,
(	88016	)	,
(	87904	)	,
(	87793	)	,
(	87682	)	,
(	87572	)	,
(	87462	)	,
(	87352	)	,
(	87242	)	,
(	87132	)	,
(	87023	)	,
(	86914	)	,
(	86806	)	,
(	86697	)	,
(	86589	)	,
(	86481	)	,
(	86374	)	,
(	86266	)	,
(	86159	)	,
(	86053	)	,
(	85946	)	,
(	85840	)	,
(	85734	)	,
(	85628	)	,
(	85523	)	,
(	85418	)	,
(	85313	)	,
(	85208	)	,
(	85103	)	,
(	84999	)	,
(	84895	)	,
(	84792	)	,
(	84688	)	,
(	84585	)	,
(	84482	)	,
(	84380	)	,
(	84277	)	,
(	84175	)	,
(	84073	)	,
(	83972	)	,
(	83870	)	,
(	83769	)	,
(	83668	)	,
(	83567	)	,
(	83467	)	,
(	83367	)	,
(	83267	)	,
(	83167	)	,
(	83068	)	,
(	82968	)	,
(	82869	)	,
(	82770	)	,
(	82672	)	,
(	82574	)	,
(	82476	)	,
(	82378	)	,
(	82280	)	,
(	82183	)	,
(	82086	)	,
(	81989	)	,
(	81892	)	,
(	81796	)	,
(	81699	)	,
(	81603	)	,
(	81508	)	,
(	81412	)	,
(	81317	)	,
(	81222	)	,
(	81127	)	,
(	81032	)	,
(	80938	)	,
(	80843	)	,
(	80749	)	,
(	80656	)	,
(	80562	)	,
(	80469	)	,
(	80376	)	,
(	80283	)	,
(	80190	)	,
(	80097	)	,
(	80005	)	,
(	79913	)	,
(	79821	)	,
(	79730	)	,
(	79638	)	,
(	79547	)	,
(	79456	)	,
(	79365	)	,
(	79274	)	,
(	79184	)	,
(	79094	)	,
(	79004	)	,
(	78914	)	,
(	78825	)	,
(	78735	)	,
(	78646	)	,
(	78557	)	,
(	78468	)	,
(	78380	)	,
(	78291	)	,
(	78203	)	,
(	78115	)	,
(	78027	)	,
(	77940	)	,
(	77853	)	,
(	77765	)	,
(	77678	)	,
(	77592	)	,
(	77505	)	,
(	77419	)	,
(	77332	)	,
(	77246	)	,
(	77160	)	,
(	77075	)	,
(	76989	)	,
(	76904	)	,
(	76819	)	,
(	76734	)	,
(	76649	)	,
(	76565	)	,
(	76481	)	,
(	76397	)	,
(	76313	)	,
(	76229	)	,
(	76145	)	,
(	76062	)	,
(	75979	)	,
(	75896	)	,
(	75813	)	,
(	75730	)	,
(	75648	)	,
(	75565	)	,
(	75483	)	,
(	75401	)	,
(	75319	)	,
(	75238	)	,
(	75156	)	,
(	75075	)	,
(	74994	)	,
(	74913	)	,
(	74832	)	,
(	74752	)	,
(	74671	)	,
(	74591	)	,
(	74511	)	,
(	74431	)	,
(	74352	)	,
(	74272	)	,
(	74193	)	,
(	74114	)	,
(	74035	)	,
(	73956	)	,
(	73877	)	,
(	73799	)	,
(	73720	)	,
(	73642	)	,
(	73564	)	,
(	73486	)	,
(	73409	)	,
(	73331	)	,
(	73254	)	,
(	73176	)	,
(	73099	)	,
(	73023	)	,
(	72946	)	,
(	72869	)	,
(	72793	)	,
(	72717	)	,
(	72641	)	,
(	72565	)	,
(	72489	)	,
(	72413	)	,
(	72338	)	,
(	72263	)	,
(	72188	)	,
(	72113	)	,
(	72038	)	,
(	71963	)	,
(	71889	)	,
(	71814	)	,
(	71740	)	,
(	71666	)	,
(	71592	)	,
(	71518	)	,
(	71445	)	,
(	71371	)	,
(	71298	)	,
(	71225	)	,
(	71152	)	,
(	71079	)	,
(	71007	)	,
(	70934	)	,
(	70862	)	,
(	70789	)	,
(	70717	)	,
(	70645	)	,
(	70574	)	,
(	70502	)	,
(	70430	)	,
(	70359	)	,
(	70288	)	,
(	70217	)	,
(	70146	)	,
(	70075	)	,
(	70004	)	,
(	69934	)	,
(	69864	)	,
(	69793	)	,
(	69723	)	,
(	69653	)	,
(	69584	)	,
(	69514	)	,
(	69444	)	,
(	69375	)	,
(	69306	)	,
(	69237	)	,
(	69168	)	,
(	69099	)	,
(	69030	)	,
(	68962	)	,
(	68893	)	,
(	68825	)	,
(	68757	)	,
(	68689	)	,
(	68621	)	,
(	68553	)	,
(	68486	)	,
(	68418	)	,
(	68351	)	,
(	68284	)	,
(	68217	)	,
(	68150	)	,
(	68083	)	,
(	68016	)	,
(	67950	)	,
(	67883	)	,
(	67817	)	,
(	67751	)	,
(	67685	)	,
(	67619	)	,
(	67553	)	,
(	67487	)	,
(	67422	)	,
(	67356	)	,
(	67291	)	,
(	67226	)	,
(	67161	)	,
(	67096	)	,
(	67031	)	,
(	66967	)	,
(	66902	)	,
(	66838	)	,
(	66774	)	,
(	66709	)	,
(	66645	)	,
(	66581	)	,
(	66518	)	,
(	66454	)	,
(	66390	)	,
(	66327	)	,
(	66264	)	,
(	66201	)	,
(	66138	)	,
(	66075	)	,
(	66012	)	,
(	65949	)	,
(	65887	)	,
(	65824	)	,
(	65762	)	,
(	65700	)	,
(	65637	)	,
(	65575	)	,
(	65514	)	,
(	65452	)	,
(	65390	)	,
(	65329	)	,
(	65267	)	,
(	65206	)	,
(	65145	)	,
(	65084	)	,
(	65023	)	,
(	64962	)	,
(	64901	)	,
(	64841	)	,
(	64780	)	,
(	64720	)	,
(	64660	)	,
(	64599	)	,
(	64539	)	,
(	64480	)	,
(	64420	)	,
(	64360	)	,
(	64300	)	,
(	64241	)	,
(	64182	)	,
(	64122	)	,
(	64063	)	,
(	64004	)	,
(	63945	)	,
(	63886	)	,
(	63828	)	,
(	63769	)	,
(	63710	)	,
(	63652	)	,
(	63594	)	,
(	63536	)	,
(	63478	)	,
(	63420	)	,
(	63362	)	,
(	63304	)	,
(	63246	)	,
(	63189	)	,
(	63131	)	,
(	63074	)	,
(	63017	)	,
(	62960	)	,
(	62903	)	,
(	62846	)	,
(	62789	)	,
(	62732	)	,
(	62675	)	,
(	62619	)	,
(	62563	)	,
(	62506	)	,
(	62450	)	,
(	62394	)	,
(	62338	)	,
(	62282	)	,
(	62226	)	,
(	62170	)	,
(	62115	)	,
(	62059	)	,
(	62004	)	,
(	61949	)	,
(	61893	)	,
(	61838	)	,
(	61783	)	,
(	61728	)	,
(	61674	)	,
(	61619	)	,
(	61564	)	,
(	61510	)	,
(	61455	)	,
(	61401	)	,
(	61347	)	,
(	61293	)	,
(	61238	)	,
(	61185	)	,
(	61131	)	,
(	61077	)	,
(	61023	)	,
(	60970	)	,
(	60916	)	,
(	60863	)	,
(	60809	)	,
(	60756	)	,
(	60703	)	,
(	60650	)	,
(	60597	)	,
(	60544	)	,
(	60492	)	,
(	60439	)	,
(	60386	)	,
(	60334	)	,
(	60282	)	,
(	60229	)	,
(	60177	)	,
(	60125	)	,
(	60073	)	,
(	60021	)	,
(	59969	)	,
(	59918	)	,
(	59866	)	,
(	59814	)	,
(	59763	)	,
(	59711	)	,
(	59660	)	,
(	59609	)	,
(	59558	)	,
(	59507	)	,
(	59456	)	,
(	59405	)	,
(	59354	)	,
(	59304	)	,
(	59253	)	,
(	59202	)	,
(	59152	)	,
(	59102	)	,
(	59051	)	,
(	59001	)	,
(	58951	)	,
(	58901	)	,
(	58851	)	,
(	58801	)	,
(	58752	)	,
(	58702	)	,
(	58652	)	,
(	58603	)	,
(	58553	)	,
(	58504	)	,
(	58455	)	,
(	58406	)	,
(	58357	)	,
(	58308	)	,
(	58259	)	,
(	58210	)	,
(	58161	)	,
(	58113	)	,
(	58064	)	,
(	58015	)	,
(	57967	)	,
(	57919	)	,
(	57870	)	,
(	57822	)	,
(	57774	)	,
(	57726	)	,
(	57678	)	,
(	57630	)	,
(	57582	)	,
(	57535	)	,
(	57487	)	,
(	57440	)	,
(	57392	)	,
(	57345	)	,
(	57297	)	,
(	57250	)	,
(	57203	)	,
(	57156	)	,
(	57109	)	,
(	57062	)	,
(	57015	)	,
(	56968	)	,
(	56922	)	,
(	56875	)	,
(	56829	)	,
(	56782	)	,
(	56736	)	,
(	56689	)	,
(	56643	)	,
(	56597	)	,
(	56551	)	,
(	56505	)	,
(	56459	)	,
(	56413	)	,
(	56367	)	,
(	56322	)	,
(	56276	)	,
(	56230	)	,
(	56185	)	,
(	56139	)	,
(	56094	)	,
(	56049	)	,
(	56004	)	,
(	55958	)	,
(	55913	)	,
(	55868	)	,
(	55824	)	,
(	55779	)	,
(	55734	)	,
(	55689	)	,
(	55645	)	,
(	55600	)	,
(	55556	)	,
(	55511	)	,
(	55467	)	,
(	55423	)	,
(	55378	)	,
(	55334	)	,
(	55290	)	,
(	55246	)	,
(	55202	)	,
(	55158	)	,
(	55115	)	,
(	55071	)	,
(	55027	)	,
(	54984	)	,
(	54940	)	,
(	54897	)	,
(	54853	)	,
(	54810	)	,
(	54767	)	,
(	54724	)	,
(	54681	)	,
(	54638	)	,
(	54595	)	,
(	54552	)	,
(	54509	)	,
(	54466	)	,
(	54424	)	,
(	54381	)	,
(	54338	)	,
(	54296	)	,
(	54253	)	,
(	54211	)	,
(	54169	)	,
(	54127	)	,
(	54084	)	,
(	54042	)	,
(	54000	)	,
(	53958	)	,
(	53916	)	,
(	53875	)	,
(	53833	)	,
(	53791	)	,
(	53750	)	,
(	53708	)	,
(	53666	)	,
(	53625	)	,
(	53584	)	,
(	53542	)	,
(	53501	)	,
(	53460	)	,
(	53419	)	,
(	53378	)	,
(	53337	)	,
(	53296	)	,
(	53255	)	,
(	53214	)	,
(	53173	)	,
(	53133	)	,
(	53092	)	,
(	53052	)	,
(	53011	)	,
(	52971	)	,
(	52930	)	,
(	52890	)	,
(	52850	)	,
(	52809	)	,
(	52769	)	,
(	52729	)	,
(	52689	)	,
(	52649	)	,
(	52609	)	,
(	52570	)	,
(	52530	)	,
(	52490	)	,
(	52450	)	,
(	52411	)	,
(	52371	)	,
(	52332	)	,
(	52293	)	,
(	52253	)	,
(	52214	)	,
(	52175	)	,
(	52135	)	,
(	52096	)	,
(	52057	)	,
(	52018	)	,
(	51979	)	,
(	51940	)	,
(	51902	)	,
(	51863	)	,
(	51824	)	,
(	51786	)	,
(	51747	)	,
(	51708	)	,
(	51670	)	,
(	51632	)	,
(	51593	)	,
(	51555	)	,
(	51517	)	,
(	51478	)	,
(	51440	)	,
(	51402	)	,
(	51364	)	,
(	51326	)	,
(	51288	)	,
(	51251	)	,
(	51213	)	,
(	51175	)	,
(	51137	)	,
(	51100	)	,
(	51062	)	,
(	51025	)	,
(	50987	)	,
(	50950	)	,
(	50912	)	,
(	50875	)	,
(	50838	)	,
(	50801	)	,
(	50763	)	,
(	50726	)	,
(	50689	)	,
(	50652	)	,
(	50615	)	,
(	50579	)	,
(	50542	)	,
(	50505	)	,
(	50468	)	,
(	50432	)	,
(	50395	)	,
(	50359	)	,
(	50322	)	,
(	50286	)	,
(	50249	)	,
(	50213	)	,
(	50177	)	,
(	50140	)	,
(	50104	)	,
(	50068	)	,
(	50032	)	,
(	49996	)	,
(	49960	)	,
(	49924	)	,
(	49888	)	,
(	49852	)	,
(	49817	)	,
(	49781	)	,
(	49745	)	,
(	49710	)	,
(	49674	)	,
(	49639	)	,
(	49603	)	,
(	49568	)	,
(	49532	)	,
(	49497	)	,
(	49462	)	,
(	49427	)	,
(	49391	)	,
(	49356	)	,
(	49321	)	,
(	49286	)	,
(	49251	)	,
(	49216	)	,
(	49182	)	,
(	49147	)	,
(	49112	)	,
(	49077	)	,
(	49043	)	,
(	49008	)	,
(	48974	)	,
(	48939	)	,
(	48905	)	,
(	48870	)	,
(	48836	)	,
(	48801	)	,
(	48767	)	,
(	48733	)	,
(	48699	)	,
(	48665	)	,
(	48631	)	,
(	48597	)	,
(	48563	)	,
(	48529	)	,
(	48495	)	,
(	48461	)	,
(	48427	)	,
(	48393	)	,
(	48360	)	,
(	48326	)	,
(	48292	)	,
(	48259	)	,
(	48225	)	,
(	48192	)	,
(	48158	)	,
(	48125	)	,
(	48092	)	,
(	48058	)	,
(	48025	)	,
(	47992	)	,
(	47959	)	,
(	47926	)	,
(	47893	)	,
(	47860	)	,
(	47827	)	,
(	47794	)	,
(	47761	)	,
(	47728	)	,
(	47695	)	,
(	47663	)	,
(	47630	)	,
(	47597	)	,
(	47565	)	,
(	47532	)	,
(	47500	)	,
(	47467	)	,
(	47435	)	,
(	47402	)	,
(	47370	)	,
(	47338	)	,
(	47305	)	,
(	47273	)	,
(	47241	)	,
(	47209	)	,
(	47177	)	,
(	47145	)	,
(	47113	)	,
(	47081	)	,
(	47049	)	,
(	47017	)	,
(	46985	)	,
(	46954	)	,
(	46922	)	,
(	46890	)	,
(	46859	)	,
(	46827	)	,
(	46795	)	,
(	46764	)	,
(	46732	)	,
(	46701	)	,
(	46670	)	,
(	46638	)	,
(	46607	)	,
(	46576	)	,
(	46545	)	,
(	46513	)	,
(	46482	)	,
(	46451	)	,
(	46420	)	,
(	46389	)	,
(	46358	)	,
(	46327	)	,
(	46296	)	,
(	46265	)	,
(	46235	)	,
(	46204	)	,
(	46173	)	,
(	46142	)	,
(	46112	)	,
(	46081	)	,
(	46051	)	,
(	46020	)	,
(	45990	)	,
(	45959	)	,
(	45929	)	,
(	45899	)	,
(	45868	)	,
(	45838	)	,
(	45808	)	,
(	45777	)	,
(	45747	)	,
(	45717	)	,
(	45687	)	,
(	45657	)	,
(	45627	)	,
(	45597	)	,
(	45567	)	,
(	45537	)	,
(	45507	)	,
(	45478	)	,
(	45448	)	,
(	45418	)	,
(	45389	)	,
(	45359	)	,
(	45329	)	,
(	45300	)	,
(	45270	)	,
(	45241	)	,
(	45211	)	,
(	45182	)	,
(	45152	)	,
(	45123	)	,
(	45094	)	,
(	45065	)	,
(	45035	)	,
(	45006	)	,
(	44977	)	,
(	44948	)	,
(	44919	)	,
(	44890	)	,
(	44861	)	,
(	44832	)	,
(	44803	)	,
(	44774	)	,
(	44745	)	,
(	44716	)	,
(	44688	)	,
(	44659	)	,
(	44630	)	,
(	44601	)	,
(	44573	)	,
(	44544	)	,
(	44516	)	,
(	44487	)	,
(	44459	)	,
(	44430	)	,
(	44402	)	,
(	44373	)	,
(	44345	)	,
(	44317	)	,
(	44289	)	,
(	44260	)	,
(	44232	)	,
(	44204	)	,
(	44176	)	,
(	44148	)	,
(	44120	)	,
(	44092	)	,
(	44064	)	,
(	44036	)	,
(	44008	)	,
(	43980	)	,
(	43952	)	,
(	43924	)	,
(	43897	)	,
(	43869	)	,
(	43841	)	,
(	43814	)	,
(	43786	)	,
(	43758	)	,
(	43731	)	,
(	43703	)	,
(	43676	)	,
(	43648	)	,
(	43621	)	,
(	43593	)	,
(	43566	)	,
(	43539	)	,
(	43512	)	,
(	43484	)	,
(	43457	)	,
(	43430	)	,
(	43403	)	,
(	43376	)	,
(	43349	)	,
(	43322	)	,
(	43295	)	,
(	43268	)	,
(	43241	)	,
(	43214	)	,
(	43187	)	,
(	43160	)	,
(	43133	)	,
(	43106	)	,
(	43080	)	,
(	43053	)	,
(	43026	)	,
(	43000	)	,
(	42973	)	,
(	42946	)	,
(	42920	)	,
(	42893	)	,
(	42867	)	,
(	42840	)	,
(	42814	)	,
(	42788	)	,
(	42761	)	,
(	42735	)	,
(	42709	)	,
(	42683	)	,
(	42656	)	,
(	42630	)	,
(	42604	)	,
(	42578	)	,
(	42552	)	,
(	42526	)	,
(	42500	)	,
(	42474	)	,
(	42448	)	,
(	42422	)	,
(	42396	)	,
(	42370	)	,
(	42344	)	,
(	42318	)	,
(	42293	)	,
(	42267	)	,
(	42241	)	,
(	42215	)	,
(	42190	)	,
(	42164	)	,
(	42139	)	,
(	42113	)	,
(	42088	)	,
(	42062	)	,
(	42037	)	,
(	42011	)	,
(	41986	)	,
(	41960	)	,
(	41935	)	,
(	41910	)	,
(	41884	)	,
(	41859	)	,
(	41834	)	,
(	41809	)	,
(	41784	)	,
(	41759	)	,
(	41733	)	,
(	41708	)	,
(	41683	)	,
(	41658	)	,
(	41633	)	,
(	41608	)	,
(	41583	)	,
(	41559	)	,
(	41534	)	,
(	41509	)	,
(	41484	)	,
(	41459	)	,
(	41435	)	,
(	41410	)	,
(	41385	)	,
(	41361	)	,
(	41336	)	,
(	41311	)	,
(	41287	)	,
(	41262	)	,
(	41238	)	,
(	41213	)	,
(	41189	)	,
(	41164	)	,
(	41140	)	,
(	41116	)	,
(	41091	)	,
(	41067	)	,
(	41043	)	,
(	41019	)	,
(	40994	)	,
(	40970	)	,
(	40946	)	,
(	40922	)	,
(	40898	)	,
(	40874	)	,
(	40850	)	,
(	40826	)	,
(	40802	)	,
(	40778	)	,
(	40754	)	,
(	40730	)	,
(	40706	)	,
(	40682	)	,
(	40658	)	,
(	40635	)	,
(	40611	)	,
(	40587	)	,
(	40563	)	,
(	40540	)	,
(	40516	)	,
(	40492	)	,
(	40469	)	,
(	40445	)	,
(	40422	)	,
(	40398	)	,
(	40375	)	,
(	40351	)	,
(	40328	)	,
(	40304	)	,
(	40281	)	,
(	40258	)	,
(	40234	)	,
(	40211	)	,
(	40188	)	,
(	40165	)	,
(	40141	)	,
(	40118	)	,
(	40095	)	,
(	40072	)	,
(	40049	)	,
(	40026	)	,
(	40003	)	,
(	39980	)	,
(	39957	)	,
(	39934	)	,
(	39911	)	,
(	39888	)	,
(	39865	)	,
(	39842	)	,
(	39819	)	,
(	39796	)	,
(	39773	)	,
(	39751	)	,
(	39728	)	,
(	39705	)	,
(	39683	)	,
(	39660	)	,
(	39637	)	,
(	39615	)	,
(	39592	)	,
(	39569	)	,
(	39547	)	,
(	39524	)	,
(	39502	)	,
(	39480	)	,
(	39457	)	,
(	39435	)	,
(	39412	)	,
(	39390	)	,
(	39368	)	,
(	39345	)	,
(	39323	)	,
(	39301	)	,
(	39279	)	,
(	39256	)	,
(	39234	)	,
(	39212	)	,
(	39190	)	,
(	39168	)	,
(	39146	)	,
(	39124	)	,
(	39102	)	,
(	39080	)	,
(	39058	)	,
(	39036	)	,
(	39014	)	,
(	38992	)	,
(	38970	)	,
(	38948	)	,
(	38926	)	,
(	38904	)	,
(	38883	)	,
(	38861	)	,
(	38839	)	,
(	38817	)	,
(	38796	)	,
(	38774	)	,
(	38752	)	,
(	38731	)	,
(	38709	)	,
(	38688	)	,
(	38666	)	,
(	38645	)	,
(	38623	)	,
(	38602	)	,
(	38580	)	,
(	38559	)	,
(	38537	)	,
(	38516	)	,
(	38495	)	,
(	38473	)	,
(	38452	)	,
(	38431	)	,
(	38410	)	,
(	38388	)	,
(	38367	)	,
(	38346	)	,
(	38325	)	,
(	38304	)	,
(	38282	)	,
(	38261	)	,
(	38240	)	,
(	38219	)	,
(	38198	)	,
(	38177	)	,
(	38156	)	,
(	38135	)	,
(	38114	)	,
(	38093	)	,
(	38073	)	,
(	38052	)	,
(	38031	)	,
(	38010	)	,
(	37989	)	,
(	37969	)	,
(	37948	)	,
(	37927	)	,
(	37906	)	,
(	37886	)	,
(	37865	)	,
(	37844	)	,
(	37824	)	,
(	37803	)	,
(	37783	)	,
(	37762	)	,
(	37742	)	,
(	37721	)	,
(	37701	)	,
(	37680	)	,
(	37660	)	,
(	37639	)	,
(	37619	)	,
(	37599	)	,
(	37578	)	,
(	37558	)	,
(	37538	)	,
(	37517	)	,
(	37497	)	,
(	37477	)	,
(	37457	)	,
(	37436	)	,
(	37416	)	,
(	37396	)	,
(	37376	)	,
(	37356	)	,
(	37336	)	,
(	37316	)	,
(	37296	)	,
(	37276	)	,
(	37256	)	,
(	37236	)	,
(	37216	)	,
(	37196	)	,
(	37176	)	,
(	37156	)	,
(	37136	)	,
(	37116	)	,
(	37096	)	,
(	37077	)	,
(	37057	)	,
(	37037	)	,
(	37017	)	,
(	36998	)	,
(	36978	)	,
(	36958	)	,
(	36939	)	,
(	36919	)	,
(	36899	)	,
(	36880	)	,
(	36860	)	,
(	36841	)	,
(	36821	)	,
(	36802	)	,
(	36782	)	,
(	36763	)	,
(	36743	)	,
(	36724	)	,
(	36704	)	,
(	36685	)	,
(	36665	)	,
(	36646	)	,
(	36627	)	,
(	36608	)	,
(	36588	)	,
(	36569	)	,
(	36550	)	,
(	36530	)	,
(	36511	)	,
(	36492	)	,
(	36473	)	,
(	36454	)	,
(	36435	)	,
(	36416	)	,
(	36396	)	,
(	36377	)	,
(	36358	)	,
(	36339	)	,
(	36320	)	,
(	36301	)	,
(	36282	)	,
(	36263	)	,
(	36244	)	,
(	36226	)	,
(	36207	)	,
(	36188	)	,
(	36169	)	,
(	36150	)	,
(	36131	)	,
(	36113	)	,
(	36094	)	,
(	36075	)	,
(	36056	)	,
(	36038	)	,
(	36019	)	,
(	36000	)	,
(	35982	)	,
(	35963	)	,
(	35944	)	,
(	35926	)	,
(	35907	)	,
(	35889	)	,
(	35870	)	,
(	35852	)	,
(	35833	)	,
(	35815	)	,
(	35796	)	,
(	35778	)	,
(	35759	)	,
(	35741	)	,
(	35722	)	,
(	35704	)	,
(	35686	)	,
(	35667	)	,
(	35649	)	,
(	35631	)	,
(	35613	)	,
(	35594	)	,
(	35576	)	,
(	35558	)	,
(	35540	)	,
(	35521	)	,
(	35503	)	,
(	35485	)	,
(	35467	)	,
(	35449	)	,
(	35431	)	,
(	35413	)	,
(	35395	)	,
(	35377	)	,
(	35359	)	,
(	35341	)	,
(	35323	)	,
(	35305	)	,
(	35287	)	,
(	35269	)	,
(	35251	)	,
(	35233	)	,
(	35215	)	,
(	35197	)	,
(	35180	)	,
(	35162	)	,
(	35144	)	,
(	35126	)	,
(	35108	)	,
(	35091	)	,
(	35073	)	,
(	35055	)	,
(	35038	)	,
(	35020	)	,
(	35002	)	,
(	34985	)	,
(	34967	)	,
(	34949	)	,
(	34932	)	,
(	34914	)	,
(	34897	)	,
(	34879	)	,
(	34862	)	,
(	34844	)	,
(	34827	)	,
(	34809	)	,
(	34792	)	,
(	34774	)	,
(	34757	)	,
(	34740	)	,
(	34722	)	,
(	34705	)	,
(	34688	)	,
(	34670	)	,
(	34653	)	,
(	34636	)	,
(	34618	)	,
(	34601	)	,
(	34584	)	,
(	34567	)	,
(	34549	)	,
(	34532	)	,
(	34515	)	,
(	34498	)	,
(	34481	)	,
(	34464	)	,
(	34447	)	,
(	34430	)	,
(	34413	)	,
(	34395	)	,
(	34378	)	,
(	34361	)	,
(	34344	)	,
(	34327	)	,
(	34310	)	,
(	34294	)	,
(	34277	)	,
(	34260	)	,
(	34243	)	,
(	34226	)	,
(	34209	)	,
(	34192	)	,
(	34175	)	,
(	34159	)	,
(	34142	)	,
(	34125	)	,
(	34108	)	,
(	34092	)	,
(	34075	)	,
(	34058	)	,
(	34041	)	,
(	34025	)	,
(	34008	)	,
(	33991	)	,
(	33975	)	,
(	33958	)	,
(	33942	)	,
(	33925	)	,
(	33908	)	,
(	33892	)	,
(	33875	)	,
(	33859	)	,
(	33842	)	,
(	33826	)	,
(	33809	)	,
(	33793	)	,
(	33776	)	,
(	33760	)	,
(	33744	)	,
(	33727	)	,
(	33711	)	,
(	33695	)	,
(	33678	)	,
(	33662	)	,
(	33646	)	,
(	33629	)	,
(	33613	)	,
(	33597	)	,
(	33580	)	,
(	33564	)	,
(	33548	)	,
(	33532	)	,
(	33516	)	,
(	33499	)	,
(	33483	)	,
(	33467	)	,
(	33451	)	,
(	33435	)	,
(	33419	)	,
(	33403	)	,
(	33387	)	,
(	33371	)	,
(	33355	)	,
(	33339	)	,
(	33323	)	,
(	33307	)	,
(	33291	)	,
(	33275	)	,
(	33259	)	,
(	33243	)	,
(	33227	)	,
(	33211	)	,
(	33195	)	,
(	33179	)	,
(	33164	)	,
(	33148	)	,
(	33132	)	,
(	33116	)	,
(	33100	)	,
(	33085	)	,
(	33069	)	,
(	33053	)	,
(	33037	)	,
(	33022	)	,
(	33006	)	,
(	32990	)	,
(	32975	)	,
(	32959	)	,
(	32943	)	,
(	32928	)	,
(	32912	)	,
(	32896	)	,
(	32881	)	,
(	32865	)	,
(	32850	)	,
(	32834	)	,
(	32819	)	,
(	32803	)	,
(	32788	)	,
(	32772	)	,
(	32757	)	,
(	32741	)	,
(	32726	)	,
(	32711	)	,
(	32695	)	,
(	32680	)	,
(	32664	)	,
(	32649	)	,
(	32634	)	,
(	32618	)	,
(	32603	)	,
(	32588	)	,
(	32572	)	,
(	32557	)	,
(	32542	)	,
(	32527	)	,
(	32511	)	,
(	32496	)	,
(	32481	)	,
(	32466	)	,
(	32451	)	,
(	32436	)	,
(	32420	)	,
(	32405	)	,
(	32390	)	,
(	32375	)	,
(	32360	)	,
(	32345	)	,
(	32330	)	,
(	32315	)	,
(	32300	)	,
(	32285	)	,
(	32270	)	,
(	32255	)	,
(	32240	)	,
(	32225	)	,
(	32210	)	,
(	32195	)	,
(	32180	)	,
(	32165	)	,
(	32150	)	,
(	32135	)	,
(	32120	)	,
(	32106	)	,
(	32091	)	,
(	32076	)	,
(	32061	)	,
(	32046	)	,
(	32032	)	,
(	32017	)	,
(	32002	)	,
(	31987	)	,
(	31973	)	,
(	31958	)	,
(	31943	)	,
(	31928	)	,
(	31914	)	,
(	31899	)	,
(	31885	)	,
(	31870	)	,
(	31855	)	,
(	31841	)	,
(	31826	)	,
(	31811	)	,
(	31797	)	,
(	31782	)	,
(	31768	)	,
(	31753	)	,
(	31739	)	,
(	31724	)	,
(	31710	)	,
(	31695	)	,
(	31681	)	,
(	31666	)	,
(	31652	)	,
(	31638	)	,
(	31623	)	,
(	31609	)	,
(	31594	)	,
(	31580	)	,
(	31566	)	,
(	31551	)	,
(	31537	)	,
(	31523	)	,
(	31508	)	,
(	31494	)	,
(	31480	)	,
(	31466	)	,
(	31451	)	,
(	31437	)	,
(	31423	)	,
(	31409	)	,
(	31394	)	,
(	31380	)	,
(	31366	)	,
(	31352	)	,
(	31338	)	,
(	31324	)	,
(	31309	)	,
(	31295	)	,
(	31281	)	,
(	31267	)	,
(	31253	)	,
(	31239	)	,
(	31225	)	,
(	31211	)	,
(	31197	)	,
(	31183	)	,
(	31169	)	,
(	31155	)	,
(	31141	)	,
(	31127	)	,
(	31113	)	,
(	31099	)	,
(	31085	)	,
(	31071	)	,
(	31057	)	,
(	31044	)	,
(	31030	)	,
(	31016	)	,
(	31002	)	,
(	30988	)	,
(	30974	)	,
(	30961	)	,
(	30947	)	,
(	30933	)	,
(	30919	)	,
(	30905	)	,
(	30892	)	,
(	30878	)	,
(	30864	)	,
(	30850	)	,
(	30837	)	,
(	30823	)	,
(	30809	)	,
(	30796	)	,
(	30782	)	,
(	30768	)	,
(	30755	)	,
(	30741	)	,
(	30728	)	,
(	30714	)	,
(	30700	)	,
(	30687	)	,
(	30673	)	,
(	30660	)	,
(	30646	)	,
(	30633	)	,
(	30619	)	,
(	30606	)	,
(	30592	)	,
(	30579	)	,
(	30565	)	,
(	30552	)	,
(	30538	)	,
(	30525	)	,
(	30512	)	,
(	30498	)	,
(	30485	)	,
(	30471	)	,
(	30458	)	,
(	30445	)	,
(	30431	)	,
(	30418	)	,
(	30405	)	,
(	30391	)	,
(	30378	)	,
(	30365	)	,
(	30352	)	,
(	30338	)	,
(	30325	)	,
(	30312	)	,
(	30299	)	,
(	30285	)	,
(	30272	)	,
(	30259	)	,
(	30246	)	,
(	30233	)	,
(	30220	)	,
(	30206	)	,
(	30193	)	,
(	30180	)	,
(	30167	)	,
(	30154	)	,
(	30141	)	,
(	30128	)	,
(	30115	)	,
(	30102	)	,
(	30089	)	,
(	30076	)	,
(	30063	)	,
(	30050	)	,
(	30037	)	,
(	30024	)	,
(	30011	)	,
(	29998	)	,
(	29985	)	,
(	29972	)	,
(	29959	)	,
(	29946	)	,
(	29933	)	,
(	29920	)	,
(	29907	)	,
(	29894	)	,
(	29881	)	,
(	29869	)	,
(	29856	)	,
(	29843	)	,
(	29830	)	,
(	29817	)	,
(	29804	)	,
(	29792	)	,
(	29779	)	,
(	29766	)	,
(	29753	)	,
(	29741	)	,
(	29728	)	,
(	29715	)	,
(	29702	)	,
(	29690	)	,
(	29677	)	,
(	29664	)	,
(	29652	)	,
(	29639	)	,
(	29626	)	,
(	29614	)	,
(	29601	)	,
(	29589	)	,
(	29576	)	,
(	29563	)	,
(	29551	)	,
(	29538	)	,
(	29526	)	,
(	29513	)	,
(	29501	)	,
(	29488	)	,
(	29476	)	,
(	29463	)	,
(	29451	)	,
(	29438	)	,
(	29426	)	,
(	29413	)	,
(	29401	)	,
(	29388	)	,
(	29376	)	,
(	29363	)	,
(	29351	)	,
(	29339	)	,
(	29326	)	,
(	29314	)	,
(	29301	)	,
(	29289	)	,
(	29277	)	,
(	29264	)	,
(	29252	)	,
(	29240	)	,
(	29227	)	,
(	29215	)	,
(	29203	)	,
(	29191	)	,
(	29178	)	,
(	29166	)	,
(	29154	)	,
(	29142	)	,
(	29129	)	,
(	29117	)	,
(	29105	)	,
(	29093	)	,
(	29081	)	,
(	29068	)	,
(	29056	)	,
(	29044	)	,
(	29032	)	,
(	29020	)	,
(	29008	)	,
(	28996	)	,
(	28983	)	,
(	28971	)	,
(	28959	)	,
(	28947	)	,
(	28935	)	,
(	28923	)	,
(	28911	)	,
(	28899	)	,
(	28887	)	,
(	28875	)	,
(	28863	)	,
(	28851	)	,
(	28839	)	,
(	28827	)	,
(	28815	)	,
(	28803	)	,
(	28791	)	,
(	28779	)	,
(	28767	)	,
(	28755	)	,
(	28744	)	,
(	28732	)	,
(	28720	)	,
(	28708	)	,
(	28696	)	,
(	28684	)	,
(	28672	)	,
(	28661	)	,
(	28649	)	,
(	28637	)	,
(	28625	)	,
(	28613	)	,
(	28602	)	,
(	28590	)	,
(	28578	)	,
(	28566	)	,
(	28554	)	,
(	28543	)	,
(	28531	)	,
(	28519	)	,
(	28508	)	,
(	28496	)	,
(	28484	)	,
(	28473	)	,
(	28461	)	,
(	28449	)	,
(	28438	)	,
(	28426	)	,
(	28414	)	,
(	28403	)	,
(	28391	)	,
(	28379	)	,
(	28368	)	,
(	28356	)	,
(	28345	)	,
(	28333	)	,
(	28322	)	,
(	28310	)	,
(	28298	)	,
(	28287	)	,
(	28275	)	,
(	28264	)	,
(	28252	)	,
(	28241	)	,
(	28229	)	,
(	28218	)	,
(	28207	)	,
(	28195	)	,
(	28184	)	,
(	28172	)	,
(	28161	)	,
(	28149	)	,
(	28138	)	,
(	28127	)	,
(	28115	)	,
(	28104	)	,
(	28092	)	,
(	28081	)	,
(	28070	)	,
(	28058	)	,
(	28047	)	,
(	28036	)	,
(	28024	)	,
(	28013	)	,
(	28002	)	,
(	27991	)	,
(	27979	)	,
(	27968	)	,
(	27957	)	,
(	27945	)	,
(	27934	)	,
(	27923	)	,
(	27912	)	,
(	27901	)	,
(	27889	)	,
(	27878	)	,
(	27867	)	,
(	27856	)	,
(	27845	)	,
(	27833	)	,
(	27822	)	,
(	27811	)	,
(	27800	)	,
(	27789	)	,
(	27778	)	,
(	27767	)	,
(	27756	)	,
(	27744	)	,
(	27733	)	,
(	27722	)	,
(	27711	)	,
(	27700	)	,
(	27689	)	,
(	27678	)	,
(	27667	)	,
(	27656	)	,
(	27645	)	,
(	27634	)	,
(	27623	)	,
(	27612	)	,
(	27601	)	,
(	27590	)	,
(	27579	)	,
(	27568	)	,
(	27557	)	,
(	27546	)	,
(	27535	)	,
(	27525	)	,
(	27514	)	,
(	27503	)	,
(	27492	)	,
(	27481	)	,
(	27470	)	,
(	27459	)	,
(	27448	)	,
(	27438	)	,
(	27427	)	,
(	27416	)	,
(	27405	)	,
(	27394	)	,
(	27383	)	,
(	27373	)	,
(	27362	)	,
(	27351	)	,
(	27340	)	,
(	27330	)	,
(	27319	)	,
(	27308	)	,
(	27297	)	,
(	27287	)	,
(	27276	)	,
(	27265	)	,
(	27254	)	,
(	27244	)	,
(	27233	)	,
(	27222	)	,
(	27212	)	,
(	27201	)	,
(	27190	)	,
(	27180	)	,
(	27169	)	,
(	27159	)	,
(	27148	)	,
(	27137	)	,
(	27127	)	,
(	27116	)	,
(	27106	)	,
(	27095	)	,
(	27084	)	,
(	27074	)	,
(	27063	)	,
(	27053	)	,
(	27042	)	,
(	27032	)	,
(	27021	)	,
(	27011	)	,
(	27000	)	,
(	26990	)	,
(	26979	)	,
(	26969	)	,
(	26958	)	,
(	26948	)	,
(	26937	)	,
(	26927	)	,
(	26916	)	,
(	26906	)	,
(	26896	)	,
(	26885	)	,
(	26875	)	,
(	26864	)	,
(	26854	)	,
(	26844	)	,
(	26833	)	,
(	26823	)	,
(	26813	)	,
(	26802	)	,
(	26792	)	,
(	26782	)	,
(	26771	)	,
(	26761	)	,
(	26751	)	,
(	26740	)	,
(	26730	)	,
(	26720	)	,
(	26709	)	,
(	26699	)	,
(	26689	)	,
(	26679	)	,
(	26668	)	,
(	26658	)	,
(	26648	)	,
(	26638	)	,
(	26627	)	,
(	26617	)	,
(	26607	)	,
(	26597	)	,
(	26587	)	,
(	26577	)	,
(	26566	)	,
(	26556	)	,
(	26546	)	,
(	26536	)	,
(	26526	)	,
(	26516	)	,
(	26506	)	,
(	26495	)	,
(	26485	)	,
(	26475	)	,
(	26465	)	,
(	26455	)	,
(	26445	)	,
(	26435	)	,
(	26425	)	,
(	26415	)	,
(	26405	)	,
(	26395	)	,
(	26385	)	,
(	26375	)	,
(	26365	)	,
(	26355	)	,
(	26345	)	,
(	26335	)	,
(	26325	)	,
(	26315	)	,
(	26305	)	,
(	26295	)	,
(	26285	)	,
(	26275	)	,
(	26265	)	,
(	26255	)	,
(	26245	)	,
(	26235	)	,
(	26225	)	,
(	26215	)	,
(	26205	)	,
(	26196	)	,
(	26186	)	,
(	26176	)	,
(	26166	)	,
(	26156	)	,
(	26146	)	,
(	26136	)	,
(	26127	)	,
(	26117	)	,
(	26107	)	,
(	26097	)	,
(	26087	)	,
(	26078	)	,
(	26068	)	,
(	26058	)	,
(	26048	)	,
(	26038	)	,
(	26029	)	,
(	26019	)	,
(	26009	)	,
(	25999	)	,
(	25990	)	,
(	25980	)	,
(	25970	)	,
(	25961	)	,
(	25951	)	,
(	25941	)	,
(	25931	)	,
(	25922	)	,
(	25912	)	,
(	25902	)	,
(	25893	)	,
(	25883	)	,
(	25873	)	,
(	25864	)	,
(	25854	)	,
(	25845	)	,
(	25835	)	,
(	25825	)	,
(	25816	)	,
(	25806	)	,
(	25797	)	,
(	25787	)	,
(	25777	)	,
(	25768	)	,
(	25758	)	,
(	25749	)	,
(	25739	)	,
(	25730	)	,
(	25720	)	,
(	25711	)	,
(	25701	)	,
(	25692	)	,
(	25682	)	,
(	25673	)	,
(	25663	)	,
(	25654	)	,
(	25644	)	,
(	25635	)	,
(	25625	)	,
(	25616	)	,
(	25606	)	,
(	25597	)	,
(	25587	)	,
(	25578	)	,
(	25569	)	,
(	25559	)	,
(	25550	)	,
(	25540	)	,
(	25531	)	,
(	25522	)	,
(	25512	)	,
(	25503	)	,
(	25494	)	,
(	25484	)	,
(	25475	)	,
(	25466	)	,
(	25456	)	,
(	25447	)	,
(	25438	)	,
(	25428	)	,
(	25419	)	,
(	25410	)	,
(	25400	)	,
(	25391	)	,
(	25382	)	,
(	25372	)	,
(	25363	)	,
(	25354	)	,
(	25345	)	,
(	25335	)	,
(	25326	)	,
(	25317	)	,
(	25308	)	,
(	25299	)	,
(	25289	)	,
(	25280	)	,
(	25271	)	,
(	25262	)	,
(	25253	)	,
(	25243	)	,
(	25234	)	,
(	25225	)	,
(	25216	)	,
(	25207	)	,
(	25198	)	,
(	25188	)	,
(	25179	)	,
(	25170	)	,
(	25161	)	,
(	25152	)	,
(	25143	)	,
(	25134	)	,
(	25125	)	,
(	25116	)	,
(	25106	)	,
(	25097	)	,
(	25088	)	,
(	25079	)	,
(	25070	)	,
(	25061	)	,
(	25052	)	,
(	25043	)	,
(	25034	)	,
(	25025	)	,
(	25016	)	,
(	25007	)	,
(	24998	)	,
(	24989	)	,
(	24980	)	,
(	24971	)	,
(	24962	)	,
(	24953	)	,
(	24944	)	,
(	24935	)	,
(	24926	)	,
(	24917	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)	,
(	250000	)


);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	
	yeet : process(index)
	begin
		if(index < 0) then
			Divisor <= 250000;
		elsif (index > 4095) then
			Divisor <= 250000;
		else
			Divisor <= Divisors(index);
		end if;
	end process;
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
