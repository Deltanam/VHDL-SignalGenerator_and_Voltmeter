
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY BuzzAmp_Lookup IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      index      	 :  IN    integer;                           
      Amplitude     :  OUT   STD_LOGIC_VECTOR(11 DOWNTO 0)
		);
END BuzzAmp_Lookup;

ARCHITECTURE behavior OF BuzzAmp_Lookup IS

type array_1d is array (0 to 4095) of integer;

constant BuzzAmps : array_1d := (				
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4	)	,
(	6	)	,
(	7	)	,
(	9	)	,
(	10	)	,
(	12	)	,
(	13	)	,
(	15	)	,
(	16	)	,
(	18	)	,
(	19	)	,
(	21	)	,
(	22	)	,
(	24	)	,
(	25	)	,
(	27	)	,
(	28	)	,
(	30	)	,
(	31	)	,
(	33	)	,
(	34	)	,
(	36	)	,
(	37	)	,
(	39	)	,
(	40	)	,
(	42	)	,
(	43	)	,
(	45	)	,
(	46	)	,
(	48	)	,
(	49	)	,
(	51	)	,
(	52	)	,
(	54	)	,
(	55	)	,
(	57	)	,
(	58	)	,
(	60	)	,
(	61	)	,
(	63	)	,
(	64	)	,
(	66	)	,
(	67	)	,
(	69	)	,
(	70	)	,
(	72	)	,
(	73	)	,
(	75	)	,
(	76	)	,
(	78	)	,
(	79	)	,
(	81	)	,
(	82	)	,
(	84	)	,
(	85	)	,
(	87	)	,
(	88	)	,
(	90	)	,
(	91	)	,
(	93	)	,
(	94	)	,
(	96	)	,
(	97	)	,
(	99	)	,
(	100	)	,
(	102	)	,
(	103	)	,
(	105	)	,
(	106	)	,
(	108	)	,
(	109	)	,
(	111	)	,
(	112	)	,
(	114	)	,
(	115	)	,
(	117	)	,
(	118	)	,
(	120	)	,
(	121	)	,
(	123	)	,
(	124	)	,
(	126	)	,
(	127	)	,
(	129	)	,
(	130	)	,
(	132	)	,
(	133	)	,
(	135	)	,
(	136	)	,
(	138	)	,
(	139	)	,
(	141	)	,
(	142	)	,
(	144	)	,
(	145	)	,
(	147	)	,
(	148	)	,
(	150	)	,
(	151	)	,
(	153	)	,
(	154	)	,
(	156	)	,
(	157	)	,
(	159	)	,
(	160	)	,
(	162	)	,
(	163	)	,
(	165	)	,
(	166	)	,
(	168	)	,
(	169	)	,
(	171	)	,
(	172	)	,
(	174	)	,
(	175	)	,
(	177	)	,
(	178	)	,
(	180	)	,
(	181	)	,
(	183	)	,
(	184	)	,
(	186	)	,
(	187	)	,
(	189	)	,
(	190	)	,
(	192	)	,
(	193	)	,
(	195	)	,
(	196	)	,
(	198	)	,
(	199	)	,
(	201	)	,
(	202	)	,
(	204	)	,
(	205	)	,
(	207	)	,
(	208	)	,
(	210	)	,
(	211	)	,
(	213	)	,
(	214	)	,
(	216	)	,
(	217	)	,
(	219	)	,
(	220	)	,
(	222	)	,
(	223	)	,
(	225	)	,
(	226	)	,
(	228	)	,
(	229	)	,
(	231	)	,
(	232	)	,
(	234	)	,
(	235	)	,
(	237	)	,
(	238	)	,
(	240	)	,
(	241	)	,
(	243	)	,
(	244	)	,
(	245	)	,
(	247	)	,
(	248	)	,
(	250	)	,
(	251	)	,
(	253	)	,
(	254	)	,
(	256	)	,
(	257	)	,
(	259	)	,
(	260	)	,
(	262	)	,
(	263	)	,
(	265	)	,
(	266	)	,
(	268	)	,
(	269	)	,
(	271	)	,
(	272	)	,
(	274	)	,
(	275	)	,
(	277	)	,
(	278	)	,
(	280	)	,
(	281	)	,
(	283	)	,
(	284	)	,
(	286	)	,
(	287	)	,
(	289	)	,
(	290	)	,
(	292	)	,
(	293	)	,
(	295	)	,
(	296	)	,
(	298	)	,
(	299	)	,
(	301	)	,
(	302	)	,
(	304	)	,
(	305	)	,
(	307	)	,
(	308	)	,
(	310	)	,
(	311	)	,
(	313	)	,
(	314	)	,
(	316	)	,
(	317	)	,
(	319	)	,
(	320	)	,
(	322	)	,
(	323	)	,
(	325	)	,
(	326	)	,
(	328	)	,
(	329	)	,
(	331	)	,
(	332	)	,
(	334	)	,
(	335	)	,
(	337	)	,
(	338	)	,
(	340	)	,
(	341	)	,
(	343	)	,
(	344	)	,
(	346	)	,
(	347	)	,
(	349	)	,
(	350	)	,
(	352	)	,
(	353	)	,
(	355	)	,
(	356	)	,
(	358	)	,
(	359	)	,
(	361	)	,
(	362	)	,
(	364	)	,
(	365	)	,
(	367	)	,
(	368	)	,
(	370	)	,
(	371	)	,
(	373	)	,
(	374	)	,
(	376	)	,
(	377	)	,
(	379	)	,
(	380	)	,
(	382	)	,
(	383	)	,
(	385	)	,
(	386	)	,
(	388	)	,
(	389	)	,
(	391	)	,
(	392	)	,
(	394	)	,
(	395	)	,
(	397	)	,
(	398	)	,
(	400	)	,
(	401	)	,
(	403	)	,
(	404	)	,
(	406	)	,
(	407	)	,
(	409	)	,
(	410	)	,
(	412	)	,
(	413	)	,
(	415	)	,
(	416	)	,
(	418	)	,
(	419	)	,
(	421	)	,
(	422	)	,
(	424	)	,
(	425	)	,
(	427	)	,
(	428	)	,
(	430	)	,
(	431	)	,
(	433	)	,
(	434	)	,
(	436	)	,
(	437	)	,
(	439	)	,
(	440	)	,
(	442	)	,
(	443	)	,
(	445	)	,
(	446	)	,
(	448	)	,
(	449	)	,
(	451	)	,
(	452	)	,
(	454	)	,
(	455	)	,
(	457	)	,
(	458	)	,
(	460	)	,
(	461	)	,
(	463	)	,
(	464	)	,
(	466	)	,
(	467	)	,
(	469	)	,
(	470	)	,
(	472	)	,
(	473	)	,
(	475	)	,
(	476	)	,
(	478	)	,
(	479	)	,
(	481	)	,
(	482	)	,
(	484	)	,
(	485	)	,
(	486	)	,
(	488	)	,
(	489	)	,
(	491	)	,
(	492	)	,
(	494	)	,
(	495	)	,
(	497	)	,
(	498	)	,
(	500	)	,
(	501	)	,
(	503	)	,
(	504	)	,
(	506	)	,
(	507	)	,
(	509	)	,
(	510	)	,
(	512	)	,
(	513	)	,
(	515	)	,
(	516	)	,
(	518	)	,
(	519	)	,
(	521	)	,
(	522	)	,
(	524	)	,
(	525	)	,
(	527	)	,
(	528	)	,
(	530	)	,
(	531	)	,
(	533	)	,
(	534	)	,
(	536	)	,
(	537	)	,
(	539	)	,
(	540	)	,
(	542	)	,
(	543	)	,
(	545	)	,
(	546	)	,
(	548	)	,
(	549	)	,
(	551	)	,
(	552	)	,
(	554	)	,
(	555	)	,
(	557	)	,
(	558	)	,
(	560	)	,
(	561	)	,
(	563	)	,
(	564	)	,
(	566	)	,
(	567	)	,
(	569	)	,
(	570	)	,
(	572	)	,
(	573	)	,
(	575	)	,
(	576	)	,
(	578	)	,
(	579	)	,
(	581	)	,
(	582	)	,
(	584	)	,
(	585	)	,
(	587	)	,
(	588	)	,
(	590	)	,
(	591	)	,
(	593	)	,
(	594	)	,
(	596	)	,
(	597	)	,
(	599	)	,
(	600	)	,
(	602	)	,
(	603	)	,
(	605	)	,
(	606	)	,
(	608	)	,
(	609	)	,
(	611	)	,
(	612	)	,
(	614	)	,
(	615	)	,
(	617	)	,
(	618	)	,
(	620	)	,
(	621	)	,
(	623	)	,
(	624	)	,
(	626	)	,
(	627	)	,
(	629	)	,
(	630	)	,
(	632	)	,
(	633	)	,
(	635	)	,
(	636	)	,
(	638	)	,
(	639	)	,
(	641	)	,
(	642	)	,
(	644	)	,
(	645	)	,
(	647	)	,
(	648	)	,
(	650	)	,
(	651	)	,
(	653	)	,
(	654	)	,
(	656	)	,
(	657	)	,
(	659	)	,
(	660	)	,
(	662	)	,
(	663	)	,
(	665	)	,
(	666	)	,
(	668	)	,
(	669	)	,
(	671	)	,
(	672	)	,
(	674	)	,
(	675	)	,
(	677	)	,
(	678	)	,
(	680	)	,
(	681	)	,
(	683	)	,
(	684	)	,
(	686	)	,
(	687	)	,
(	689	)	,
(	690	)	,
(	692	)	,
(	693	)	,
(	695	)	,
(	696	)	,
(	698	)	,
(	699	)	,
(	701	)	,
(	702	)	,
(	704	)	,
(	705	)	,
(	707	)	,
(	708	)	,
(	710	)	,
(	711	)	,
(	713	)	,
(	714	)	,
(	716	)	,
(	717	)	,
(	719	)	,
(	720	)	,
(	722	)	,
(	723	)	,
(	725	)	,
(	726	)	,
(	727	)	,
(	729	)	,
(	730	)	,
(	732	)	,
(	733	)	,
(	735	)	,
(	736	)	,
(	738	)	,
(	739	)	,
(	741	)	,
(	742	)	,
(	744	)	,
(	745	)	,
(	747	)	,
(	748	)	,
(	750	)	,
(	751	)	,
(	753	)	,
(	754	)	,
(	756	)	,
(	757	)	,
(	759	)	,
(	760	)	,
(	762	)	,
(	763	)	,
(	765	)	,
(	766	)	,
(	768	)	,
(	769	)	,
(	771	)	,
(	772	)	,
(	774	)	,
(	775	)	,
(	777	)	,
(	778	)	,
(	780	)	,
(	781	)	,
(	783	)	,
(	784	)	,
(	786	)	,
(	787	)	,
(	789	)	,
(	790	)	,
(	792	)	,
(	793	)	,
(	795	)	,
(	796	)	,
(	798	)	,
(	799	)	,
(	801	)	,
(	802	)	,
(	804	)	,
(	805	)	,
(	807	)	,
(	808	)	,
(	810	)	,
(	811	)	,
(	813	)	,
(	814	)	,
(	816	)	,
(	817	)	,
(	819	)	,
(	820	)	,
(	822	)	,
(	823	)	,
(	825	)	,
(	826	)	,
(	828	)	,
(	829	)	,
(	831	)	,
(	832	)	,
(	834	)	,
(	835	)	,
(	837	)	,
(	838	)	,
(	840	)	,
(	841	)	,
(	843	)	,
(	844	)	,
(	846	)	,
(	847	)	,
(	849	)	,
(	850	)	,
(	852	)	,
(	853	)	,
(	855	)	,
(	856	)	,
(	858	)	,
(	859	)	,
(	861	)	,
(	862	)	,
(	864	)	,
(	865	)	,
(	867	)	,
(	868	)	,
(	870	)	,
(	871	)	,
(	873	)	,
(	874	)	,
(	876	)	,
(	877	)	,
(	879	)	,
(	880	)	,
(	882	)	,
(	883	)	,
(	885	)	,
(	886	)	,
(	888	)	,
(	889	)	,
(	891	)	,
(	892	)	,
(	894	)	,
(	895	)	,
(	897	)	,
(	898	)	,
(	900	)	,
(	901	)	,
(	903	)	,
(	904	)	,
(	906	)	,
(	907	)	,
(	909	)	,
(	910	)	,
(	912	)	,
(	913	)	,
(	915	)	,
(	916	)	,
(	918	)	,
(	919	)	,
(	921	)	,
(	922	)	,
(	924	)	,
(	925	)	,
(	927	)	,
(	928	)	,
(	930	)	,
(	931	)	,
(	933	)	,
(	934	)	,
(	936	)	,
(	937	)	,
(	939	)	,
(	940	)	,
(	942	)	,
(	943	)	,
(	945	)	,
(	946	)	,
(	948	)	,
(	949	)	,
(	951	)	,
(	952	)	,
(	954	)	,
(	955	)	,
(	957	)	,
(	958	)	,
(	960	)	,
(	961	)	,
(	963	)	,
(	964	)	,
(	966	)	,
(	967	)	,
(	968	)	,
(	970	)	,
(	971	)	,
(	973	)	,
(	974	)	,
(	976	)	,
(	977	)	,
(	979	)	,
(	980	)	,
(	982	)	,
(	983	)	,
(	985	)	,
(	986	)	,
(	988	)	,
(	989	)	,
(	991	)	,
(	992	)	,
(	994	)	,
(	995	)	,
(	997	)	,
(	998	)	,
(	1000	)	,
(	1001	)	,
(	1003	)	,
(	1004	)	,
(	1006	)	,
(	1007	)	,
(	1009	)	,
(	1010	)	,
(	1012	)	,
(	1013	)	,
(	1015	)	,
(	1016	)	,
(	1018	)	,
(	1019	)	,
(	1021	)	,
(	1022	)	,
(	1024	)	,
(	1025	)	,
(	1027	)	,
(	1028	)	,
(	1030	)	,
(	1031	)	,
(	1033	)	,
(	1034	)	,
(	1036	)	,
(	1037	)	,
(	1039	)	,
(	1040	)	,
(	1042	)	,
(	1043	)	,
(	1045	)	,
(	1046	)	,
(	1048	)	,
(	1049	)	,
(	1051	)	,
(	1052	)	,
(	1054	)	,
(	1055	)	,
(	1057	)	,
(	1058	)	,
(	1060	)	,
(	1061	)	,
(	1063	)	,
(	1064	)	,
(	1066	)	,
(	1067	)	,
(	1069	)	,
(	1070	)	,
(	1072	)	,
(	1073	)	,
(	1075	)	,
(	1076	)	,
(	1078	)	,
(	1079	)	,
(	1081	)	,
(	1082	)	,
(	1084	)	,
(	1085	)	,
(	1087	)	,
(	1088	)	,
(	1090	)	,
(	1091	)	,
(	1093	)	,
(	1094	)	,
(	1096	)	,
(	1097	)	,
(	1099	)	,
(	1100	)	,
(	1102	)	,
(	1103	)	,
(	1105	)	,
(	1106	)	,
(	1108	)	,
(	1109	)	,
(	1111	)	,
(	1112	)	,
(	1114	)	,
(	1115	)	,
(	1117	)	,
(	1118	)	,
(	1120	)	,
(	1121	)	,
(	1123	)	,
(	1124	)	,
(	1126	)	,
(	1127	)	,
(	1129	)	,
(	1130	)	,
(	1132	)	,
(	1133	)	,
(	1135	)	,
(	1136	)	,
(	1138	)	,
(	1139	)	,
(	1141	)	,
(	1142	)	,
(	1144	)	,
(	1145	)	,
(	1147	)	,
(	1148	)	,
(	1150	)	,
(	1151	)	,
(	1153	)	,
(	1154	)	,
(	1156	)	,
(	1157	)	,
(	1159	)	,
(	1160	)	,
(	1162	)	,
(	1163	)	,
(	1165	)	,
(	1166	)	,
(	1168	)	,
(	1169	)	,
(	1171	)	,
(	1172	)	,
(	1174	)	,
(	1175	)	,
(	1177	)	,
(	1178	)	,
(	1180	)	,
(	1181	)	,
(	1183	)	,
(	1184	)	,
(	1186	)	,
(	1187	)	,
(	1189	)	,
(	1190	)	,
(	1192	)	,
(	1193	)	,
(	1195	)	,
(	1196	)	,
(	1198	)	,
(	1199	)	,
(	1201	)	,
(	1202	)	,
(	1204	)	,
(	1205	)	,
(	1207	)	,
(	1208	)	,
(	1209	)	,
(	1211	)	,
(	1212	)	,
(	1214	)	,
(	1215	)	,
(	1217	)	,
(	1218	)	,
(	1220	)	,
(	1221	)	,
(	1223	)	,
(	1224	)	,
(	1226	)	,
(	1227	)	,
(	1229	)	,
(	1230	)	,
(	1232	)	,
(	1233	)	,
(	1235	)	,
(	1236	)	,
(	1238	)	,
(	1239	)	,
(	1241	)	,
(	1242	)	,
(	1244	)	,
(	1245	)	,
(	1247	)	,
(	1248	)	,
(	1250	)	,
(	1251	)	,
(	1253	)	,
(	1254	)	,
(	1256	)	,
(	1257	)	,
(	1259	)	,
(	1260	)	,
(	1262	)	,
(	1263	)	,
(	1265	)	,
(	1266	)	,
(	1268	)	,
(	1269	)	,
(	1271	)	,
(	1272	)	,
(	1274	)	,
(	1275	)	,
(	1277	)	,
(	1278	)	,
(	1280	)	,
(	1281	)	,
(	1283	)	,
(	1284	)	,
(	1286	)	,
(	1287	)	,
(	1289	)	,
(	1290	)	,
(	1292	)	,
(	1293	)	,
(	1295	)	,
(	1296	)	,
(	1298	)	,
(	1299	)	,
(	1301	)	,
(	1302	)	,
(	1304	)	,
(	1305	)	,
(	1307	)	,
(	1308	)	,
(	1310	)	,
(	1311	)	,
(	1313	)	,
(	1314	)	,
(	1316	)	,
(	1317	)	,
(	1319	)	,
(	1320	)	,
(	1322	)	,
(	1323	)	,
(	1325	)	,
(	1326	)	,
(	1328	)	,
(	1329	)	,
(	1331	)	,
(	1332	)	,
(	1334	)	,
(	1335	)	,
(	1337	)	,
(	1338	)	,
(	1340	)	,
(	1341	)	,
(	1343	)	,
(	1344	)	,
(	1346	)	,
(	1347	)	,
(	1349	)	,
(	1350	)	,
(	1352	)	,
(	1353	)	,
(	1355	)	,
(	1356	)	,
(	1358	)	,
(	1359	)	,
(	1361	)	,
(	1362	)	,
(	1364	)	,
(	1365	)	,
(	1367	)	,
(	1368	)	,
(	1370	)	,
(	1371	)	,
(	1373	)	,
(	1374	)	,
(	1376	)	,
(	1377	)	,
(	1379	)	,
(	1380	)	,
(	1382	)	,
(	1383	)	,
(	1385	)	,
(	1386	)	,
(	1388	)	,
(	1389	)	,
(	1391	)	,
(	1392	)	,
(	1394	)	,
(	1395	)	,
(	1397	)	,
(	1398	)	,
(	1400	)	,
(	1401	)	,
(	1403	)	,
(	1404	)	,
(	1406	)	,
(	1407	)	,
(	1409	)	,
(	1410	)	,
(	1412	)	,
(	1413	)	,
(	1415	)	,
(	1416	)	,
(	1418	)	,
(	1419	)	,
(	1421	)	,
(	1422	)	,
(	1424	)	,
(	1425	)	,
(	1427	)	,
(	1428	)	,
(	1430	)	,
(	1431	)	,
(	1433	)	,
(	1434	)	,
(	1436	)	,
(	1437	)	,
(	1439	)	,
(	1440	)	,
(	1442	)	,
(	1443	)	,
(	1445	)	,
(	1446	)	,
(	1448	)	,
(	1449	)	,
(	1451	)	,
(	1452	)	,
(	1453	)	,
(	1455	)	,
(	1456	)	,
(	1458	)	,
(	1459	)	,
(	1461	)	,
(	1462	)	,
(	1464	)	,
(	1465	)	,
(	1467	)	,
(	1468	)	,
(	1470	)	,
(	1471	)	,
(	1473	)	,
(	1474	)	,
(	1476	)	,
(	1477	)	,
(	1479	)	,
(	1480	)	,
(	1482	)	,
(	1483	)	,
(	1485	)	,
(	1486	)	,
(	1488	)	,
(	1489	)	,
(	1491	)	,
(	1492	)	,
(	1494	)	,
(	1495	)	,
(	1497	)	,
(	1498	)	,
(	1500	)	,
(	1501	)	,
(	1503	)	,
(	1504	)	,
(	1506	)	,
(	1507	)	,
(	1509	)	,
(	1510	)	,
(	1512	)	,
(	1513	)	,
(	1515	)	,
(	1516	)	,
(	1518	)	,
(	1519	)	,
(	1521	)	,
(	1522	)	,
(	1524	)	,
(	1525	)	,
(	1527	)	,
(	1528	)	,
(	1530	)	,
(	1531	)	,
(	1533	)	,
(	1534	)	,
(	1536	)	,
(	1537	)	,
(	1539	)	,
(	1540	)	,
(	1542	)	,
(	1543	)	,
(	1545	)	,
(	1546	)	,
(	1548	)	,
(	1549	)	,
(	1551	)	,
(	1552	)	,
(	1554	)	,
(	1555	)	,
(	1557	)	,
(	1558	)	,
(	1560	)	,
(	1561	)	,
(	1563	)	,
(	1564	)	,
(	1566	)	,
(	1567	)	,
(	1569	)	,
(	1570	)	,
(	1572	)	,
(	1573	)	,
(	1575	)	,
(	1576	)	,
(	1578	)	,
(	1579	)	,
(	1581	)	,
(	1582	)	,
(	1584	)	,
(	1585	)	,
(	1587	)	,
(	1588	)	,
(	1590	)	,
(	1591	)	,
(	1593	)	,
(	1594	)	,
(	1596	)	,
(	1597	)	,
(	1599	)	,
(	1600	)	,
(	1602	)	,
(	1603	)	,
(	1605	)	,
(	1606	)	,
(	1608	)	,
(	1609	)	,
(	1611	)	,
(	1612	)	,
(	1614	)	,
(	1615	)	,
(	1617	)	,
(	1618	)	,
(	1620	)	,
(	1621	)	,
(	1623	)	,
(	1624	)	,
(	1626	)	,
(	1627	)	,
(	1629	)	,
(	1630	)	,
(	1632	)	,
(	1633	)	,
(	1635	)	,
(	1636	)	,
(	1638	)	,
(	1639	)	,
(	1641	)	,
(	1642	)	,
(	1644	)	,
(	1645	)	,
(	1647	)	,
(	1648	)	,
(	1650	)	,
(	1651	)	,
(	1653	)	,
(	1654	)	,
(	1656	)	,
(	1657	)	,
(	1659	)	,
(	1660	)	,
(	1662	)	,
(	1663	)	,
(	1665	)	,
(	1666	)	,
(	1668	)	,
(	1669	)	,
(	1671	)	,
(	1672	)	,
(	1674	)	,
(	1675	)	,
(	1677	)	,
(	1678	)	,
(	1680	)	,
(	1681	)	,
(	1683	)	,
(	1684	)	,
(	1686	)	,
(	1687	)	,
(	1689	)	,
(	1690	)	,
(	1692	)	,
(	1693	)	,
(	1694	)	,
(	1696	)	,
(	1697	)	,
(	1699	)	,
(	1700	)	,
(	1702	)	,
(	1703	)	,
(	1705	)	,
(	1706	)	,
(	1708	)	,
(	1709	)	,
(	1711	)	,
(	1712	)	,
(	1714	)	,
(	1715	)	,
(	1717	)	,
(	1718	)	,
(	1720	)	,
(	1721	)	,
(	1723	)	,
(	1724	)	,
(	1726	)	,
(	1727	)	,
(	1729	)	,
(	1730	)	,
(	1732	)	,
(	1733	)	,
(	1735	)	,
(	1736	)	,
(	1738	)	,
(	1739	)	,
(	1741	)	,
(	1742	)	,
(	1744	)	,
(	1745	)	,
(	1747	)	,
(	1748	)	,
(	1750	)	,
(	1751	)	,
(	1753	)	,
(	1754	)	,
(	1756	)	,
(	1757	)	,
(	1759	)	,
(	1760	)	,
(	1762	)	,
(	1763	)	,
(	1765	)	,
(	1766	)	,
(	1768	)	,
(	1769	)	,
(	1771	)	,
(	1772	)	,
(	1774	)	,
(	1775	)	,
(	1777	)	,
(	1778	)	,
(	1780	)	,
(	1781	)	,
(	1783	)	,
(	1784	)	,
(	1786	)	,
(	1787	)	,
(	1789	)	,
(	1790	)	,
(	1792	)	,
(	1793	)	,
(	1795	)	,
(	1796	)	,
(	1798	)	,
(	1799	)	,
(	1801	)	,
(	1802	)	,
(	1804	)	,
(	1805	)	,
(	1807	)	,
(	1808	)	,
(	1810	)	,
(	1811	)	,
(	1813	)	,
(	1814	)	,
(	1816	)	,
(	1817	)	,
(	1819	)	,
(	1820	)	,
(	1822	)	,
(	1823	)	,
(	1825	)	,
(	1826	)	,
(	1828	)	,
(	1829	)	,
(	1831	)	,
(	1832	)	,
(	1834	)	,
(	1835	)	,
(	1837	)	,
(	1838	)	,
(	1840	)	,
(	1841	)	,
(	1843	)	,
(	1844	)	,
(	1846	)	,
(	1847	)	,
(	1849	)	,
(	1850	)	,
(	1852	)	,
(	1853	)	,
(	1855	)	,
(	1856	)	,
(	1858	)	,
(	1859	)	,
(	1861	)	,
(	1862	)	,
(	1864	)	,
(	1865	)	,
(	1867	)	,
(	1868	)	,
(	1870	)	,
(	1871	)	,
(	1873	)	,
(	1874	)	,
(	1876	)	,
(	1877	)	,
(	1879	)	,
(	1880	)	,
(	1882	)	,
(	1883	)	,
(	1885	)	,
(	1886	)	,
(	1888	)	,
(	1889	)	,
(	1891	)	,
(	1892	)	,
(	1894	)	,
(	1895	)	,
(	1897	)	,
(	1898	)	,
(	1900	)	,
(	1901	)	,
(	1903	)	,
(	1904	)	,
(	1906	)	,
(	1907	)	,
(	1909	)	,
(	1910	)	,
(	1912	)	,
(	1913	)	,
(	1915	)	,
(	1916	)	,
(	1918	)	,
(	1919	)	,
(	1921	)	,
(	1922	)	,
(	1924	)	,
(	1925	)	,
(	1927	)	,
(	1928	)	,
(	1930	)	,
(	1931	)	,
(	1933	)	,
(	1934	)	,
(	1935	)	,
(	1937	)	,
(	1938	)	,
(	1940	)	,
(	1941	)	,
(	1943	)	,
(	1944	)	,
(	1946	)	,
(	1947	)	,
(	1949	)	,
(	1950	)	,
(	1952	)	,
(	1953	)	,
(	1955	)	,
(	1956	)	,
(	1958	)	,
(	1959	)	,
(	1961	)	,
(	1962	)	,
(	1964	)	,
(	1965	)	,
(	1967	)	,
(	1968	)	,
(	1970	)	,
(	1971	)	,
(	1973	)	,
(	1974	)	,
(	1976	)	,
(	1977	)	,
(	1979	)	,
(	1980	)	,
(	1982	)	,
(	1983	)	,
(	1985	)	,
(	1986	)	,
(	1988	)	,
(	1989	)	,
(	1991	)	,
(	1992	)	,
(	1994	)	,
(	1995	)	,
(	1997	)	,
(	1998	)	,
(	2000	)	,
(	2001	)	,
(	2003	)	,
(	2004	)	,
(	2006	)	,
(	2007	)	,
(	2009	)	,
(	2010	)	,
(	2012	)	,
(	2013	)	,
(	2015	)	,
(	2016	)	,
(	2018	)	,
(	2019	)	,
(	2021	)	,
(	2022	)	,
(	2024	)	,
(	2025	)	,
(	2027	)	,
(	2028	)	,
(	2030	)	,
(	2031	)	,
(	2033	)	,
(	2034	)	,
(	2036	)	,
(	2037	)	,
(	2039	)	,
(	2040	)	,
(	2042	)	,
(	2043	)	,
(	2045	)	,
(	2046	)	,
(	2048	)	,
(	2049	)	,
(	2051	)	,
(	2052	)	,
(	2054	)	,
(	2055	)	,
(	2057	)	,
(	2058	)	,
(	2060	)	,
(	2061	)	,
(	2063	)	,
(	2064	)	,
(	2066	)	,
(	2067	)	,
(	2069	)	,
(	2070	)	,
(	2072	)	,
(	2073	)	,
(	2075	)	,
(	2076	)	,
(	2078	)	,
(	2079	)	,
(	2081	)	,
(	2082	)	,
(	2084	)	,
(	2085	)	,
(	2087	)	,
(	2088	)	,
(	2090	)	,
(	2091	)	,
(	2093	)	,
(	2094	)	,
(	2096	)	,
(	2097	)	,
(	2099	)	,
(	2100	)	,
(	2102	)	,
(	2103	)	,
(	2105	)	,
(	2106	)	,
(	2108	)	,
(	2109	)	,
(	2111	)	,
(	2112	)	,
(	2114	)	,
(	2115	)	,
(	2117	)	,
(	2118	)	,
(	2120	)	,
(	2121	)	,
(	2123	)	,
(	2124	)	,
(	2126	)	,
(	2127	)	,
(	2129	)	,
(	2130	)	,
(	2132	)	,
(	2133	)	,
(	2135	)	,
(	2136	)	,
(	2138	)	,
(	2139	)	,
(	2141	)	,
(	2142	)	,
(	2144	)	,
(	2145	)	,
(	2147	)	,
(	2148	)	,
(	2150	)	,
(	2151	)	,
(	2153	)	,
(	2154	)	,
(	2156	)	,
(	2157	)	,
(	2159	)	,
(	2160	)	,
(	2162	)	,
(	2163	)	,
(	2165	)	,
(	2166	)	,
(	2168	)	,
(	2169	)	,
(	2171	)	,
(	2172	)	,
(	2174	)	,
(	2175	)	,
(	2176	)	,
(	2178	)	,
(	2179	)	,
(	2181	)	,
(	2182	)	,
(	2184	)	,
(	2185	)	,
(	2187	)	,
(	2188	)	,
(	2190	)	,
(	2191	)	,
(	2193	)	,
(	2194	)	,
(	2196	)	,
(	2197	)	,
(	2199	)	,
(	2200	)	,
(	2202	)	,
(	2203	)	,
(	2205	)	,
(	2206	)	,
(	2208	)	,
(	2209	)	,
(	2211	)	,
(	2212	)	,
(	2214	)	,
(	2215	)	,
(	2217	)	,
(	2218	)	,
(	2220	)	,
(	2221	)	,
(	2223	)	,
(	2224	)	,
(	2226	)	,
(	2227	)	,
(	2229	)	,
(	2230	)	,
(	2232	)	,
(	2233	)	,
(	2235	)	,
(	2236	)	,
(	2238	)	,
(	2239	)	,
(	2241	)	,
(	2242	)	,
(	2244	)	,
(	2245	)	,
(	2247	)	,
(	2248	)	,
(	2250	)	,
(	2251	)	,
(	2253	)	,
(	2254	)	,
(	2256	)	,
(	2257	)	,
(	2259	)	,
(	2260	)	,
(	2262	)	,
(	2263	)	,
(	2265	)	,
(	2266	)	,
(	2268	)	,
(	2269	)	,
(	2271	)	,
(	2272	)	,
(	2274	)	,
(	2275	)	,
(	2277	)	,
(	2278	)	,
(	2280	)	,
(	2281	)	,
(	2283	)	,
(	2284	)	,
(	2286	)	,
(	2287	)	,
(	2289	)	,
(	2290	)	,
(	2292	)	,
(	2293	)	,
(	2295	)	,
(	2296	)	,
(	2298	)	,
(	2299	)	,
(	2301	)	,
(	2302	)	,
(	2304	)	,
(	2305	)	,
(	2307	)	,
(	2308	)	,
(	2310	)	,
(	2311	)	,
(	2313	)	,
(	2314	)	,
(	2316	)	,
(	2317	)	,
(	2319	)	,
(	2320	)	,
(	2322	)	,
(	2323	)	,
(	2325	)	,
(	2326	)	,
(	2328	)	,
(	2329	)	,
(	2331	)	,
(	2332	)	,
(	2334	)	,
(	2335	)	,
(	2337	)	,
(	2338	)	,
(	2340	)	,
(	2341	)	,
(	2343	)	,
(	2344	)	,
(	2346	)	,
(	2347	)	,
(	2349	)	,
(	2350	)	,
(	2352	)	,
(	2353	)	,
(	2355	)	,
(	2356	)	,
(	2358	)	,
(	2359	)	,
(	2361	)	,
(	2362	)	,
(	2364	)	,
(	2365	)	,
(	2367	)	,
(	2368	)	,
(	2370	)	,
(	2371	)	,
(	2373	)	,
(	2374	)	,
(	2376	)	,
(	2377	)	,
(	2379	)	,
(	2380	)	,
(	2382	)	,
(	2383	)	,
(	2385	)	,
(	2386	)	,
(	2388	)	,
(	2389	)	,
(	2391	)	,
(	2392	)	,
(	2394	)	,
(	2395	)	,
(	2397	)	,
(	2398	)	,
(	2400	)	,
(	2401	)	,
(	2403	)	,
(	2404	)	,
(	2406	)	,
(	2407	)	,
(	2409	)	,
(	2410	)	,
(	2412	)	,
(	2413	)	,
(	2415	)	,
(	2416	)	,
(	2417	)	,
(	2419	)	,
(	2420	)	,
(	2422	)	,
(	2423	)	,
(	2425	)	,
(	2426	)	,
(	2428	)	,
(	2429	)	,
(	2431	)	,
(	2432	)	,
(	2434	)	,
(	2435	)	,
(	2437	)	,
(	2438	)	,
(	2440	)	,
(	2441	)	,
(	2443	)	,
(	2444	)	,
(	2446	)	,
(	2447	)	,
(	2449	)	,
(	2450	)	,
(	2452	)	,
(	2453	)	,
(	2455	)	,
(	2456	)	,
(	2458	)	,
(	2459	)	,
(	2461	)	,
(	2462	)	,
(	2464	)	,
(	2465	)	,
(	2467	)	,
(	2468	)	,
(	2470	)	,
(	2471	)	,
(	2473	)	,
(	2474	)	,
(	2476	)	,
(	2477	)	,
(	2479	)	,
(	2480	)	,
(	2482	)	,
(	2483	)	,
(	2485	)	,
(	2486	)	,
(	2488	)	,
(	2489	)	,
(	2491	)	,
(	2492	)	,
(	2494	)	,
(	2495	)	,
(	2497	)	,
(	2498	)	,
(	2500	)	,
(	2501	)	,
(	2503	)	,
(	2504	)	,
(	2506	)	,
(	2507	)	,
(	2509	)	,
(	2510	)	,
(	2512	)	,
(	2513	)	,
(	2515	)	,
(	2516	)	,
(	2518	)	,
(	2519	)	,
(	2521	)	,
(	2522	)	,
(	2524	)	,
(	2525	)	,
(	2527	)	,
(	2528	)	,
(	2530	)	,
(	2531	)	,
(	2533	)	,
(	2534	)	,
(	2536	)	,
(	2537	)	,
(	2539	)	,
(	2540	)	,
(	2542	)	,
(	2543	)	,
(	2545	)	,
(	2546	)	,
(	2548	)	,
(	2549	)	,
(	2551	)	,
(	2552	)	,
(	2554	)	,
(	2555	)	,
(	2557	)	,
(	2558	)	,
(	2560	)	,
(	2561	)	,
(	2563	)	,
(	2564	)	,
(	2566	)	,
(	2567	)	,
(	2569	)	,
(	2570	)	,
(	2572	)	,
(	2573	)	,
(	2575	)	,
(	2576	)	,
(	2578	)	,
(	2579	)	,
(	2581	)	,
(	2582	)	,
(	2584	)	,
(	2585	)	,
(	2587	)	,
(	2588	)	,
(	2590	)	,
(	2591	)	,
(	2593	)	,
(	2594	)	,
(	2596	)	,
(	2597	)	,
(	2599	)	,
(	2600	)	,
(	2602	)	,
(	2603	)	,
(	2605	)	,
(	2606	)	,
(	2608	)	,
(	2609	)	,
(	2611	)	,
(	2612	)	,
(	2614	)	,
(	2615	)	,
(	2617	)	,
(	2618	)	,
(	2620	)	,
(	2621	)	,
(	2623	)	,
(	2624	)	,
(	2626	)	,
(	2627	)	,
(	2629	)	,
(	2630	)	,
(	2632	)	,
(	2633	)	,
(	2635	)	,
(	2636	)	,
(	2638	)	,
(	2639	)	,
(	2641	)	,
(	2642	)	,
(	2644	)	,
(	2645	)	,
(	2647	)	,
(	2648	)	,
(	2650	)	,
(	2651	)	,
(	2653	)	,
(	2654	)	,
(	2656	)	,
(	2657	)	,
(	2658	)	,
(	2660	)	,
(	2661	)	,
(	2663	)	,
(	2664	)	,
(	2666	)	,
(	2667	)	,
(	2669	)	,
(	2670	)	,
(	2672	)	,
(	2673	)	,
(	2675	)	,
(	2676	)	,
(	2678	)	,
(	2679	)	,
(	2681	)	,
(	2682	)	,
(	2684	)	,
(	2685	)	,
(	2687	)	,
(	2688	)	,
(	2690	)	,
(	2691	)	,
(	2693	)	,
(	2694	)	,
(	2696	)	,
(	2697	)	,
(	2699	)	,
(	2700	)	,
(	2702	)	,
(	2703	)	,
(	2705	)	,
(	2706	)	,
(	2708	)	,
(	2709	)	,
(	2711	)	,
(	2712	)	,
(	2714	)	,
(	2715	)	,
(	2717	)	,
(	2718	)	,
(	2720	)	,
(	2721	)	,
(	2723	)	,
(	2724	)	,
(	2726	)	,
(	2727	)	,
(	2729	)	,
(	2730	)	,
(	2732	)	,
(	2733	)	,
(	2735	)	,
(	2736	)	,
(	2738	)	,
(	2739	)	,
(	2741	)	,
(	2742	)	,
(	2744	)	,
(	2745	)	,
(	2747	)	,
(	2748	)	,
(	2750	)	,
(	2751	)	,
(	2753	)	,
(	2754	)	,
(	2756	)	,
(	2757	)	,
(	2759	)	,
(	2760	)	,
(	2762	)	,
(	2763	)	,
(	2765	)	,
(	2766	)	,
(	2768	)	,
(	2769	)	,
(	2771	)	,
(	2772	)	,
(	2774	)	,
(	2775	)	,
(	2777	)	,
(	2778	)	,
(	2780	)	,
(	2781	)	,
(	2783	)	,
(	2784	)	,
(	2786	)	,
(	2787	)	,
(	2789	)	,
(	2790	)	,
(	2792	)	,
(	2793	)	,
(	2795	)	,
(	2796	)	,
(	2798	)	,
(	2799	)	,
(	2801	)	,
(	2802	)	,
(	2804	)	,
(	2805	)	,
(	2807	)	,
(	2808	)	,
(	2810	)	,
(	2811	)	,
(	2813	)	,
(	2814	)	,
(	2816	)	,
(	2817	)	,
(	2819	)	,
(	2820	)	,
(	2822	)	,
(	2823	)	,
(	2825	)	,
(	2826	)	,
(	2828	)	,
(	2829	)	,
(	2831	)	,
(	2832	)	,
(	2834	)	,
(	2835	)	,
(	2837	)	,
(	2838	)	,
(	2840	)	,
(	2841	)	,
(	2843	)	,
(	2844	)	,
(	2846	)	,
(	2847	)	,
(	2849	)	,
(	2850	)	,
(	2852	)	,
(	2853	)	,
(	2855	)	,
(	2856	)	,
(	2858	)	,
(	2859	)	,
(	2861	)	,
(	2862	)	,
(	2864	)	,
(	2865	)	,
(	2867	)	,
(	2868	)	,
(	2870	)	,
(	2871	)	,
(	2873	)	,
(	2874	)	,
(	2876	)	,
(	2877	)	,
(	2879	)	,
(	2880	)	,
(	2882	)	,
(	2883	)	,
(	2885	)	,
(	2886	)	,
(	2888	)	,
(	2889	)	,
(	2891	)	,
(	2892	)	,
(	2894	)	,
(	2895	)	,
(	2897	)	,
(	2898	)	,
(	2899	)	,
(	2901	)	,
(	2902	)	,
(	2904	)	,
(	2905	)	,
(	2907	)	,
(	2908	)	,
(	2910	)	,
(	2911	)	,
(	2913	)	,
(	2914	)	,
(	2916	)	,
(	2917	)	,
(	2919	)	,
(	2920	)	,
(	2922	)	,
(	2923	)	,
(	2925	)	,
(	2926	)	,
(	2928	)	,
(	2929	)	,
(	2931	)	,
(	2932	)	,
(	2934	)	,
(	2935	)	,
(	2937	)	,
(	2938	)	,
(	2940	)	,
(	2941	)	,
(	2943	)	,
(	2944	)	,
(	2946	)	,
(	2947	)	,
(	2949	)	,
(	2950	)	,
(	2952	)	,
(	2953	)	,
(	2955	)	,
(	2956	)	,
(	2958	)	,
(	2959	)	,
(	2961	)	,
(	2962	)	,
(	2964	)	,
(	2965	)	,
(	2967	)	,
(	2968	)	,
(	2970	)	,
(	2971	)	,
(	2973	)	,
(	2974	)	,
(	2976	)	,
(	2977	)	,
(	2979	)	,
(	2980	)	,
(	2982	)	,
(	2983	)	,
(	2985	)	,
(	2986	)	,
(	2988	)	,
(	2989	)	,
(	2991	)	,
(	2992	)	,
(	2994	)	,
(	2995	)	,
(	2997	)	,
(	2998	)	,
(	3000	)	,
(	3001	)	,
(	3003	)	,
(	3004	)	,
(	3006	)	,
(	3007	)	,
(	3009	)	,
(	3010	)	,
(	3012	)	,
(	3013	)	,
(	3015	)	,
(	3016	)	,
(	3018	)	,
(	3019	)	,
(	3021	)	,
(	3022	)	,
(	3024	)	,
(	3025	)	,
(	3027	)	,
(	3028	)	,
(	3030	)	,
(	3031	)	,
(	3033	)	,
(	3034	)	,
(	3036	)	,
(	3037	)	,
(	3039	)	,
(	3040	)	,
(	3042	)	,
(	3043	)	,
(	3045	)	,
(	3046	)	,
(	3048	)	,
(	3049	)	,
(	3051	)	,
(	3052	)	,
(	3054	)	,
(	3055	)	,
(	3057	)	,
(	3058	)	,
(	3060	)	,
(	3061	)	,
(	3063	)	,
(	3064	)	,
(	3066	)	,
(	3067	)	,
(	3069	)	,
(	3070	)	,
(	3072	)	,
(	3073	)	,
(	3075	)	,
(	3076	)	,
(	3078	)	,
(	3079	)	,
(	3081	)	,
(	3082	)	,
(	3084	)	,
(	3085	)	,
(	3087	)	,
(	3088	)	,
(	3090	)	,
(	3091	)	,
(	3093	)	,
(	3094	)	,
(	3096	)	,
(	3097	)	,
(	3099	)	,
(	3100	)	,
(	3102	)	,
(	3103	)	,
(	3105	)	,
(	3106	)	,
(	3108	)	,
(	3109	)	,
(	3111	)	,
(	3112	)	,
(	3114	)	,
(	3115	)	,
(	3117	)	,
(	3118	)	,
(	3120	)	,
(	3121	)	,
(	3123	)	,
(	3124	)	,
(	3126	)	,
(	3127	)	,
(	3129	)	,
(	3130	)	,
(	3132	)	,
(	3133	)	,
(	3135	)	,
(	3136	)	,
(	3138	)	,
(	3139	)	,
(	3141	)	,
(	3142	)	,
(	3143	)	,
(	3145	)	,
(	3146	)	,
(	3148	)	,
(	3149	)	,
(	3151	)	,
(	3152	)	,
(	3154	)	,
(	3155	)	,
(	3157	)	,
(	3158	)	,
(	3160	)	,
(	3161	)	,
(	3163	)	,
(	3164	)	,
(	3166	)	,
(	3167	)	,
(	3169	)	,
(	3170	)	,
(	3172	)	,
(	3173	)	,
(	3175	)	,
(	3176	)	,
(	3178	)	,
(	3179	)	,
(	3181	)	,
(	3182	)	,
(	3184	)	,
(	3185	)	,
(	3187	)	,
(	3188	)	,
(	3190	)	,
(	3191	)	,
(	3193	)	,
(	3194	)	,
(	3196	)	,
(	3197	)	,
(	3199	)	,
(	3200	)	,
(	3202	)	,
(	3203	)	,
(	3205	)	,
(	3206	)	,
(	3208	)	,
(	3209	)	,
(	3211	)	,
(	3212	)	,
(	3214	)	,
(	3215	)	,
(	3217	)	,
(	3218	)	,
(	3220	)	,
(	3221	)	,
(	3223	)	,
(	3224	)	,
(	3226	)	,
(	3227	)	,
(	3229	)	,
(	3230	)	,
(	3232	)	,
(	3233	)	,
(	3235	)	,
(	3236	)	,
(	3238	)	,
(	3239	)	,
(	3241	)	,
(	3242	)	,
(	3244	)	,
(	3245	)	,
(	3247	)	,
(	3248	)	,
(	3250	)	,
(	3251	)	,
(	3253	)	,
(	3254	)	,
(	3256	)	,
(	3257	)	,
(	3259	)	,
(	3260	)	,
(	3262	)	,
(	3263	)	,
(	3265	)	,
(	3266	)	,
(	3268	)	,
(	3269	)	,
(	3271	)	,
(	3272	)	,
(	3274	)	,
(	3275	)	,
(	3277	)	,
(	3278	)	,
(	3280	)	,
(	3281	)	,
(	3283	)	,
(	3284	)	,
(	3286	)	,
(	3287	)	,
(	3289	)	,
(	3290	)	,
(	3292	)	,
(	3293	)	,
(	3295	)	,
(	3296	)	,
(	3298	)	,
(	3299	)	,
(	3301	)	,
(	3302	)	,
(	3304	)	,
(	3305	)	,
(	3307	)	,
(	3308	)	,
(	3310	)	,
(	3311	)	,
(	3313	)	,
(	3314	)	,
(	3316	)	,
(	3317	)	,
(	3319	)	,
(	3320	)	,
(	3322	)	,
(	3323	)	,
(	3325	)	,
(	3326	)	,
(	3328	)	,
(	3329	)	,
(	3331	)	,
(	3332	)	,
(	3334	)	,
(	3335	)	,
(	3337	)	,
(	3338	)	,
(	3340	)	,
(	3341	)	,
(	3343	)	,
(	3344	)	,
(	3346	)	,
(	3347	)	,
(	3349	)	,
(	3350	)	,
(	3352	)	,
(	3353	)	,
(	3355	)	,
(	3356	)	,
(	3358	)	,
(	3359	)	,
(	3361	)	,
(	3362	)	,
(	3364	)	,
(	3365	)	,
(	3367	)	,
(	3368	)	,
(	3370	)	,
(	3371	)	,
(	3373	)	,
(	3374	)	,
(	3376	)	,
(	3377	)	,
(	3379	)	,
(	3380	)	,
(	3382	)	,
(	3383	)	,
(	3384	)	,
(	3386	)	,
(	3387	)	,
(	3389	)	,
(	3390	)	,
(	3392	)	,
(	3393	)	,
(	3395	)	,
(	3396	)	,
(	3398	)	,
(	3399	)	,
(	3401	)	,
(	3402	)	,
(	3404	)	,
(	3405	)	,
(	3407	)	,
(	3408	)	,
(	3410	)	,
(	3411	)	,
(	3413	)	,
(	3414	)	,
(	3416	)	,
(	3417	)	,
(	3419	)	,
(	3420	)	,
(	3422	)	,
(	3423	)	,
(	3425	)	,
(	3426	)	,
(	3428	)	,
(	3429	)	,
(	3431	)	,
(	3432	)	,
(	3434	)	,
(	3435	)	,
(	3437	)	,
(	3438	)	,
(	3440	)	,
(	3441	)	,
(	3443	)	,
(	3444	)	,
(	3446	)	,
(	3447	)	,
(	3449	)	,
(	3450	)	,
(	3452	)	,
(	3453	)	,
(	3455	)	,
(	3456	)	,
(	3458	)	,
(	3459	)	,
(	3461	)	,
(	3462	)	,
(	3464	)	,
(	3465	)	,
(	3467	)	,
(	3468	)	,
(	3470	)	,
(	3471	)	,
(	3473	)	,
(	3474	)	,
(	3476	)	,
(	3477	)	,
(	3479	)	,
(	3480	)	,
(	3482	)	,
(	3483	)	,
(	3485	)	,
(	3486	)	,
(	3488	)	,
(	3489	)	,
(	3491	)	,
(	3492	)	,
(	3494	)	,
(	3495	)	,
(	3497	)	,
(	3498	)	,
(	3500	)	,
(	3501	)	,
(	3503	)	,
(	3504	)	,
(	3506	)	,
(	3507	)	,
(	3509	)	,
(	3510	)	,
(	3512	)	,
(	3513	)	,
(	3515	)	,
(	3516	)	,
(	3518	)	,
(	3519	)	,
(	3521	)	,
(	3522	)	,
(	3524	)	,
(	3525	)	,
(	3527	)	,
(	3528	)	,
(	3530	)	,
(	3531	)	,
(	3533	)	,
(	3534	)	,
(	3536	)	,
(	3537	)	,
(	3539	)	,
(	3540	)	,
(	3542	)	,
(	3543	)	,
(	3545	)	,
(	3546	)	,
(	3548	)	,
(	3549	)	,
(	3551	)	,
(	3552	)	,
(	3554	)	,
(	3555	)	,
(	3557	)	,
(	3558	)	,
(	3560	)	,
(	3561	)	,
(	3563	)	,
(	3564	)	,
(	3566	)	,
(	3567	)	,
(	3569	)	,
(	3570	)	,
(	3572	)	,
(	3573	)	,
(	3575	)	,
(	3576	)	,
(	3578	)	,
(	3579	)	,
(	3581	)	,
(	3582	)	,
(	3584	)	,
(	3585	)	,
(	3587	)	,
(	3588	)	,
(	3590	)	,
(	3591	)	,
(	3593	)	,
(	3594	)	,
(	3596	)	,
(	3597	)	,
(	3599	)	,
(	3600	)	,
(	3602	)	,
(	3603	)	,
(	3605	)	,
(	3606	)	,
(	3608	)	,
(	3609	)	,
(	3611	)	,
(	3612	)	,
(	3614	)	,
(	3615	)	,
(	3617	)	,
(	3618	)	,
(	3620	)	,
(	3621	)	,
(	3623	)	,
(	3624	)	,
(	3625	)	,
(	3627	)	,
(	3628	)	,
(	3630	)	,
(	3631	)	,
(	3633	)	,
(	3634	)	,
(	3636	)	,
(	3637	)	,
(	3639	)	,
(	3640	)	,
(	3642	)	,
(	3643	)	,
(	3645	)	,
(	3646	)	,
(	3648	)	,
(	3649	)	,
(	3651	)	,
(	3652	)	,
(	3654	)	,
(	3655	)	,
(	3657	)	,
(	3658	)	,
(	3660	)	,
(	3661	)	,
(	3663	)	,
(	3664	)	,
(	3666	)	,
(	3667	)	,
(	3669	)	,
(	3670	)	,
(	3672	)	,
(	3673	)	,
(	3675	)	,
(	3676	)	,
(	3678	)	,
(	3679	)	,
(	3681	)	,
(	3682	)	,
(	3684	)	,
(	3685	)	,
(	3687	)	,
(	3688	)	,
(	3690	)	,
(	3691	)	,
(	3693	)	,
(	3694	)	,
(	3696	)	,
(	3697	)	,
(	3699	)	,
(	3700	)	,
(	3702	)	,
(	3703	)	,
(	3705	)	,
(	3706	)	,
(	3708	)	,
(	3709	)	,
(	3711	)	,
(	3712	)	,
(	3714	)	,
(	3715	)	,
(	3717	)	,
(	3718	)	,
(	3720	)	,
(	3721	)	,
(	3723	)	,
(	3724	)	,
(	3726	)	,
(	3727	)	,
(	3729	)	,
(	3730	)	,
(	3732	)	,
(	3733	)	,
(	3735	)	,
(	3736	)	,
(	3738	)	,
(	3739	)	,
(	3741	)	,
(	3742	)	,
(	3744	)	,
(	3745	)	,
(	3747	)	,
(	3748	)	,
(	3750	)	,
(	3751	)	,
(	3753	)	,
(	3754	)	,
(	3756	)	,
(	3757	)	,
(	3759	)	,
(	3760	)	,
(	3762	)	,
(	3763	)	,
(	3765	)	,
(	3766	)	,
(	3768	)	,
(	3769	)	,
(	3771	)	,
(	3772	)	,
(	3774	)	,
(	3775	)	,
(	3777	)	,
(	3778	)	,
(	3780	)	,
(	3781	)	,
(	3783	)	,
(	3784	)	,
(	3786	)	,
(	3787	)	,
(	3789	)	,
(	3790	)	,
(	3792	)	,
(	3793	)	,
(	3795	)	,
(	3796	)	,
(	3798	)	,
(	3799	)	,
(	3801	)	,
(	3802	)	,
(	3804	)	,
(	3805	)	,
(	3807	)	,
(	3808	)	,
(	3810	)	,
(	3811	)	,
(	3813	)	,
(	3814	)	,
(	3816	)	,
(	3817	)	,
(	3819	)	,
(	3820	)	,
(	3822	)	,
(	3823	)	,
(	3825	)	,
(	3826	)	,
(	3828	)	,
(	3829	)	,
(	3831	)	,
(	3832	)	,
(	3834	)	,
(	3835	)	,
(	3837	)	,
(	3838	)	,
(	3840	)	,
(	3841	)	,
(	3843	)	,
(	3844	)	,
(	3846	)	,
(	3847	)	,
(	3849	)	,
(	3850	)	,
(	3852	)	,
(	3853	)	,
(	3855	)	,
(	3856	)	,
(	3858	)	,
(	3859	)	,
(	3861	)	,
(	3862	)	,
(	3864	)	,
(	3865	)	,
(	3866	)	,
(	3868	)	,
(	3869	)	,
(	3871	)	,
(	3872	)	,
(	3874	)	,
(	3875	)	,
(	3877	)	,
(	3878	)	,
(	3880	)	,
(	3881	)	,
(	3883	)	,
(	3884	)	,
(	3886	)	,
(	3887	)	,
(	3889	)	,
(	3890	)	,
(	3892	)	,
(	3893	)	,
(	3895	)	,
(	3896	)	,
(	3898	)	,
(	3899	)	,
(	3901	)	,
(	3902	)	,
(	3904	)	,
(	3905	)	,
(	3907	)	,
(	3908	)	,
(	3910	)	,
(	3911	)	,
(	3913	)	,
(	3914	)	,
(	3916	)	,
(	3917	)	,
(	3919	)	,
(	3920	)	,
(	3922	)	,
(	3923	)	,
(	3925	)	,
(	3926	)	,
(	3928	)	,
(	3929	)	,
(	3931	)	,
(	3932	)	,
(	3934	)	,
(	3935	)	,
(	3937	)	,
(	3938	)	,
(	3940	)	,
(	3941	)	,
(	3943	)	,
(	3944	)	,
(	3946	)	,
(	3947	)	,
(	3949	)	,
(	3950	)	,
(	3952	)	,
(	3953	)	,
(	3955	)	,
(	3956	)	,
(	3958	)	,
(	3959	)	,
(	3961	)	,
(	3962	)	,
(	3964	)	,
(	3965	)	,
(	3967	)	,
(	3968	)	,
(	3970	)	,
(	3971	)	,
(	3973	)	,
(	3974	)	,
(	3976	)	,
(	3977	)	,
(	3979	)	,
(	3980	)	,
(	3982	)	,
(	3983	)	,
(	3985	)	,
(	3986	)	,
(	3988	)	,
(	3989	)	,
(	3991	)	,
(	3992	)	,
(	3994	)	,
(	3995	)	,
(	3997	)	,
(	3998	)	,
(	4000	)	,
(	4001	)	,
(	4003	)	,
(	4004	)	,
(	4006	)	,
(	4007	)	,
(	4009	)	,
(	4010	)	,
(	4012	)	,
(	4013	)	,
(	4015	)	,
(	4016	)	,
(	4018	)	,
(	4019	)	,
(	4021	)	,
(	4022	)	,
(	4024	)	,
(	4025	)	,
(	4027	)	,
(	4028	)	,
(	4030	)	,
(	4031	)	,
(	4033	)	,
(	4034	)	,
(	4036	)	,
(	4037	)	,
(	4039	)	,
(	4040	)	,
(	4042	)	,
(	4043	)	,
(	4045	)	,
(	4046	)	,
(	4048	)	,
(	4049	)	,
(	4051	)	,
(	4052	)	,
(	4054	)	,
(	4055	)	,
(	4057	)	,
(	4058	)	,
(	4060	)	,
(	4061	)	,
(	4063	)	,
(	4064	)	,
(	4066	)	,
(	4067	)	,
(	4069	)	,
(	4070	)	,
(	4072	)	,
(	4073	)	,
(	4075	)	,
(	4076	)	,
(	4078	)	,
(	4079	)	,
(	4081	)	,
(	4082	)	,
(	4084	)	,
(	4085	)	,
(	4087	)	,
(	4088	)	,
(	4090	)	,
(	4091	)	,
(	4093	)	,
(	4094	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)

);


begin
    -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	yeet : process(index)
	begin
		if(index < 0) then
			Amplitude <= "111111111111";
		elsif (index > 4095) then
			Amplitude <= "111111111111";
		else
			Amplitude <= std_logic_vector(to_unsigned((BuzzAmps(index)),Amplitude'length));
		end if;
	end process;
--   distance <= std_logic_vector(to_unsigned(v2d_LUTshort(to_integer(unsigned(voltage))),distance'length));
--   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
